`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
of6EBD3LINr6babdn6nrOIb1AsEkPd7G2xyAmRRNAW/kOl3oaiz8iaULce6bDa5SQjkJPIaQXORu
rA/HRghWjQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UiSveIrFN3XAU/XkbBkVqCHAe1Y8IfHlqrt1hlh346/hefiqfZ5rkZNZhu085WMw1zS47/13NO2U
IwPeYa2WCydHQxqt9PGygbmepZcU/7MwkjxkvhbcakvH3A3RrA6Gnh5K3v+/dei39oQXn2Yf9CXK
IIR/PieIVZ3eprwvjhw=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ayFi19EXsqIAV2NpuGU52JFSiOqKl1DdqYsKMX37oNaWQBp+XhZ4bdTWbpIjyl+nelyDPoK2xxQw
OVTJxJR3x0fBorId0jtI4UdxdGxSEGBx1eg6mwaxEtASxDY8AONnGRTUUfwmfuPeoQxnhjwVnpsx
JWEXyl6krJktVlxTp7k=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Vo8VffvuskbdOx6tcz3JH03fcIQMUd5iBywDqmpihLHgoPBxu/djwE2Wu7kiR88PWJaNEj7ohFZv
zvUWKDPYVlovhQo7qBUK/DuG3Pg5B2RF5Q+SWdSXKS6rhnv8wchvSPISTy1Evh4Bl+BNF+2pJpjR
un6ScX9SLQdNmBTEpFPNGZVOs/DcbJK9DBXmPSTiyHHHbfXDpfaSWm+AiLVvTRfnuAXBv/7M/M02
WIZOymomjNkDJHycP/mWLeylLBkXxUO4SkvqmQQQVgx/T8sR3FCvTDwIPiMSgDKTQVQ03RIOeFxL
orSDcWDEdOOBItv4QWWm/SrWqXlHBKJCqtkjsg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dq24mOrMj/1+5KeOJE84gP132kHy6UPWybkSrbE9jHRcQp+IWOSBgq6NFm15WNlQnrb9YRfnt75c
zPambbvh0gbhd663kLBqZtLr91IPCeVzLtiWUOBUjeSiIGUShKXR5psnKcLJzm/AlPcMuOOdAknb
qVMLbe65us8/eQ4YZvUkIQs1QQhXhBSeCKWEn+VX1I38VPPhmXaFAUr7wZ6LD+EQr7+ACsRqe4+e
KI/X+hNLEXiVP17eI6RXbvPdi6TPs/0KLYMxslkoJrxEqgC3HvQWBbIq9MjMJBvXrwajVLOcJeln
nti1B67c0vxMUqU5FFz+v43g55s+dUr1brZ+ng==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TmPPpQCnuHbpxwBtCVk229BjMiZB3o4JVmGA/AUzXfnf9eWjxDgoe99eRhNmCq+BLqtTx4PY0uC+
vnZz9Bm5W1Aip5MI6eFxOTsVZpAfzZj5GvUQXSan7jLZ7Nwr08FXPyZMi8aGJLa6EMpWHHSJGLZt
lM98SyX7y7e85kLBgh2KUdvGEL1FmKql4ryIbGABoVQw5fHgbp0Dl5d3GHGzIrDU80Isu9PmWK5O
FInWf8rU3J8RUVJbERhc68QqVlQC7ljJGHdyCVgOwJV4E8gRpvK1g7r5Ha61tO63Yf5Juk2wbFUm
BCCxeCAZSeoi6LsVj2ymtwxA/QHHUaPukwBEUw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 125824)
`protect data_block
7xLBVK/CBViFe6X3n5Pc7c9qHnK02MjfY3Pn4QClweQ6fTvddOf3qcDEK0RU3QKkHnDL5oWDilZo
PEcmv50YfLZ8+zZKo99LeBPhWvBcchgXpb0YVfPiMOzKJt4A8UIzn+nOb0PNiofKj/0/WuGJK5Nj
a8cPnHKM8OOTu38uVWU0Y08vHIKm9REIoXKCrMQ83CHHkllN6079Shp+YarfZ2YayP1w3nz3a2+X
lCCRAOuxEWhbKAVN7n7v06yroHv7PFrUiSOAoo5oPqp/2GYf7FD77yAsjqhSqaPOKDhDOgjndCQX
sRMm879+o2rmVQKmQ4QK/FxyjjXJxDWX26RcWSyhwSECqDMWdXQiBsixwOX63F2VIhpDkh9QtWhg
UfREE4+0W7p0RXRc5WKrlv9nGzP/zlgEYGaPhQN45v8jAJauw8dmDRA3ybuVPnZE6VMCa10TiucM
z8zWbXRb+Dr79BWku2juyhGnUporLHg/MiOeGjaH+eh59XtZDRzrrjZE7lscppRM+KyqJjTDXZ68
q1z5LsZ+/p9E6yXVczGx/tsP/Ix3E890vokKOZcB38fnSZMfREO0SZdm0GZ1v2ne0qo1qTueclJm
jqy2GobRH8DVFf6b7LggqThZLZTzvoWSwhcqp4UQEI/AE4cqLjd7bDjzbhhJ+ZqwPEcDS4VX/gP6
IXIuGK4W+BTqzAo8MJEYviKAepUSjaYCEDR0U/qL4pk4SMG53d5BvWBEwH4H9FT7Vd0CNbJ5P/FJ
u3V71Lt20h0ZGDmOWbEkr4rOfodQ3FzGqXpDsN6X6b919FY/iTXo08ANiBRwskp0rkd2qAUN14Gb
7VdjvLbxItG9r+Snc0qcohTnQWZYOh5rqiSWMhVw5gKBd4DWWphGesxVlEQxoQnIYCtlxiWAisZl
K1WRNP2Bxvo28RA9p56iK+kDFPk0LlHFOa9qnqU/V9S23/04z9KrRqNbxoWaH9Di5TkSry5D+LTs
QTNXwLnoOY7y3FsiiBOz0bK20XKvbUKubbM7uNvwLJRkQ5+AgVl5UJ+bjTc2A7cN2XCXFZTlsZ0z
xTf2XmEA0PbmaKA8/hJ8I9HSyonLb0b+nVhnu51iEsLvu88nfkJgIcnQCpzDPSOp2JoUUp3Gsaw1
f6ortKDH9DNCPVq/uosuOnu5gpCU7Yguojn+E7HJEa9QMuLmrM5oavu158e+p1xu2oB/E3CVrEja
cZyxbCUOXVYvPpJWS7lLeazD2kCpFU/KlcP4ALrl/aucEQPmsHzquSnqGumEGH+HJcjLI3BjrKF+
Wjlp/QExTQqltD+nHcYHEXPuRc5mpJLz6NicZstFkolBnH5hQi0Fx295lE1GCz2ZRzn2VeAOuytw
4czIkj9/TH7dYS1nwFMnHGQKjOm/mPYDwIrWsVFnYkLV1OcWJdkgSLSW3swLC5Okb53jnPt90/GL
9ycYKE+7+Y96J+3K41XhfuBQAI6HiGIFBL9fsuNJjSDGePBo0NGkLcoueTJipCOpXQi7TiRNF/Sq
/4oU8VfT0+nr/YgeRuAnnCr+BVWmORhkuiQ1sOv8vLWS3tFfqwoa21aQDx1YhDpHngUjcPZuKNIZ
zjmKLeh6GjWwU/soe//3Ir0qa/Rx/PnP9+QUhYCw8uY5d5Wp4plBgIQJUfZdjkNM9Quxmk8iAvf1
KlDXFa6H67LEs7GTVUPu3ZYjyDUe333N6diewFyCubW/ZoLb/tD2qQ1Do2o/HobHu2uQt4hM1UtZ
m3yWhIBNL4JJgfLDdSREeH16xcCjFQWoT/Le5+ijhDhEzlll6azit15PU4GAnGILKVeNSmlFfYB/
aodhUMZF5CrPC35KUir5HF/cjXD0TfuT/6uWsMGrT4MMv/tbVSiWB9LfyGn5l1TD0FJOC0MuPWQF
tC35UDrKk/m23qsK01oFGzvPaoLVscXAo+C/iyRGAQBvselFVVn5fxO9EFfMBj2xsdAsj4s2xrAX
+Y75255BqAaYy7hl1/8e18ul0KCiYTSm6LOVegPy9+G9its/pY2v/WzFLPLzgevL69owkkGqdHuI
ybW+IXVbGmWyK2eXCLLTU2iqFthKiimHg6gFtl9EGm8fYtwPD2k0mpY+cs6s2Rb5nohnQV8L3Yoe
nl0KNRwzPy1Ykj4I0eq94gcYcYGhCV8M6uPbdBWzoLLv9uN9xyNwJ87yu+HrJLQE7r+FxWTZHOzt
fNzTtKyfAS0SAraVUcW/3Dq74f8te3lre8bT5Q/4p/wQE6FWwq5POnsbuHKwtUO+7JFRFwko+qHA
5JxF8/ETfN9UksR2cgsowHInAQhC+Oz7sM002HWwEK9VThm1wRI/dTGSukigOxgClCoGL1JPqHNN
k9c7+brKHnh5LzvLItYRFEgvyTPvatTXyMUolftgQFlU3Z2ztZN377C2VpL0Li/aWzb9ftKwF/lV
aY+ee99f/SCwlYQz5bKdxbetzC1XGV0q3EvlWhW5XSrgLhDuGbPOoNpXj5GFYshmer2x79EK6B8n
LhG/EbgqR4xICsmaGjow8ZC2fGRBGtOzf1jMMLdGyLw3mKr7ZIcYryyv/v7Aiuot/aEd5QAQZuf0
E7A0XTtKWwERQRumLIjaYLSFgp+byLiTeZp0oOvVhSrgzQ7lBY7nvYDSv8r+Rt3a7zWBlguXK+JG
h+72ZZKaI4kwXAgwuS5cm6+8Ni1gWAw7A3+4bLc3Md6zWXTiHC2h7UjFTegw98Cd7++72HXW9rvx
Qpfrmxx7kxcyh+VVa4XlPM/6fpIGeSf7khhSQg8ujUZgPmVRE7SEraKATIlBAa+w3zeGj4ZKYHbK
XXPY4OgD4K4jkhLecKUJ82mjIhqhcahxBsEFiGDXA/NhRpMygWTAjtaIfJN8g+XmS5BpFxDfcmvy
lujwG/WtSBQkboOCGQoa0t82VlEfo0pix6V7aHWs/6GQWYpAbmJt1Y0or+CZhoGWDX/vPHjlmYVj
7LRpGNFri0WvjjAKoqYt9/mHfLKPJYRnyFOupjs4F5r+G2f4X0A0r7TBVHzCFqj6o7MYQ7aW0sE8
/CiFU2jY6Fda40hA2HyEW9n4C1EqY6rHKix2hLcCXR6n4A7efII+a6MWepl8Uf6OmAqcJ63tZsnK
8rynw9zagDgDeMzZBFN48DBpCoTTl9cTk5UuHX01ghwYUmM3F5abSC7nlz5gfyCLwPBfX146/yRJ
hUFDVg1lNBUffsP1e64jJMp6FpF2UzVE/lryZmlq3Wr0sgr5UxvUbI2NamSZvlo1i+GffMNdew7a
BgpMCBpkuCqgWt6q8vXrlk4oTYml6DPsOWamuwCvIqg0NPdFVFygP5JH5VUtEiZppjOqRWl9jSe/
z0xq8W7bCbszAnK1pPX1DJYwu5l1joE6WkDZUn3A65JDdabExZrthAnxlgJM0g/9J1NrJQ1MzZgq
SR/UQY5McnIbdE0ubvf1aO/zLfZlF07Wk0a4WVVQqA1fX2efnN4YPAuVMENnuTcBAIlCRU9vLWFI
ho92tATD0kvHnMBKSYeumItp+ZiJm7pB3AfC6qpeCQKXTi6nbzgLROOe8C07OgKGJJS1PxskZuND
SijvAie8YMIMDG+7ebuRfV4phGDg7u1c1ptyW9WS/7XmJD7GGN1TtJUwCWXoNdVPP/m83Sk7983S
FPAhZCQZtim91PsnOrlwAZDAY4GoKiwslWG3Lz5ZlVZ4LA7OnKq4hkf/GIJ09utWAX1uTNllqaH/
y3C7pS+oxeCaJs3r86/y/UhLaIqHdT/Bur6t4ffzchb+T08v6s5VcgZ6neGomuiwkQn7b2b/2kbz
ZXHOAk/FWS4NPqh9F2zbsNy84CcXFOjWLj9mW5KIVwdzqOvXdoyOefjj+F3CdZq074IvpE8+dhhO
M8uq5Yw18urT31YvJWDEng1qxkfb2D+C0D7ZFvuug1wGgcp2LkA7y+oQN+5RAyBEvQQsdbQeMWcE
RXbecnU+8i2oSenreIDyDJ7uVtPWprUuEuefiD1C3bKtiMYV64fPJv66K5OylMlxKem4yIn2nNnO
tqpEjzOlbmA9hYoZ1ZyUiow6nxVxS5SWRr6HaOhwsh8FeRhA0fwEWOA8ms1H1vRceXyR3w1RQIYh
bqi0U483r4Gya+5M7qdugGPDIC7a/3YAjH5CGTBIxy6quEUqwrH8NXO06jdmPW9sby/V2xlLRT6V
bi9P4b97TpJPPun7nMcex/YCTvZZeisRFejbQstqyiK/giYA3jtZDwqwJPa1Is5qJW99cJx7SybA
N843IZe4M+mobZYMIMz+DAz0Nh4LB8HCEmUyIRx1uoonai+OOgVRw6I0Qe7xE0V3YFQA8m21soX4
304wAHmN4kAHvJu5x1ceF1hHK0xv1g783Ynr1PrJXYq0cR0CIsUilUr3CWtrA616d5G/SrHoPMmM
r6+KNztOYR1CHScUFcxsrNqScXaeTX5CPLM+vwYe2/w+QvUVkQso9Qg2/FTmsaSB5Gd+bvHIdoV0
Ap2rBbFrg+VUJgJUyQPQ6rjE2Yg0xQxw+3MYGI1tj30RheBl1M5Fav/morF6okoGY9Dw+SAoYb7B
l2yv63Hw74gJy+/eL8BIfK33lPUMYTEessp6V0HCqRT2WeMma8AXG2CubN4QvqXmw1vgh7BI5ELG
4ECvYsSGxQ1GK0brBrUz+/xwFhUfEw7QjQS05P4mq7AHi2PoVOSvyXMs3/7ZcE8gIBn/vWFXh5nR
/oxlpMf+ygeR34YVyyPBh3+edKZDIYa0LZM9aXya2dDH0wfl13/KzTNBbn5TC4aOQByt3OKtYui8
ZfT/gsMDT3dyNwK1UtBuDTvHZ+msKbwdyI8+3CUV7p1IiIiJvq2shlB8daBjn7ZpH0wCgsDIpxDz
1+EfgApKRGC35+IHGoP8c4tdG2/xcTjq1abg9r5Kf2qb9eN8Ha884TdoK0FaP/yXDnZHHz5m85oY
yDB1Y3G0i7izxMgBj7h6bmnIxRgsrT7kYfJDDEafC3JUVxWsnqhbqV3TqQtKykYldqbwzfPxmaY7
2WOfwvkocwthMMmaw0xtivaemeLvt8T+xCKXz+tOuc8iWbXypRlolFeVdDl7jcpw4gRDWpeBWrFp
xudf4955l/BgcGl9hmVqUXP+W9GNT0XyphljcVUJqTKZseTTJ6ljMNII9N4I+15iVe13aiPYL8XY
dNCRB9TNeFfIsy6vwuwVvOSjwffu6hqIpQyBVUkc06ASep3RrA0fRpsxXUcLFiAe0a1MasieIXUJ
sYwOH+AEKlK9utv6WsT565gdL2TRBX4JHwMuw5tS5PaW5X2Vkmz+Kv61iryGAlhkwg6BVoB0xdUh
ATwgYbzE8WBnBbxbX7UZVuqxFwEqlKzuMx+KQXhTpgseBj4jfOHePpG7aOHksB6s9Yry09O5aosL
gjqGgWt9cs2SVrlHN2j9AvTUg0GOM42iJJCTYJ5sdLSSn7taDYm01Ibydw7Z2y4DhKNYuNYU+4XW
Tv5Kuqp/eRo0quaDJNLoh9e5uJhQ24rUOvoGv/WjVOuH3SWiF0wjLROM4qZVtIhdND/KcQXYFrjP
77kUGpSodH0I3So9Ri6D+kH+2iLFRAIE1VuNlMAvT1ISX2sjI3KFvOCXz3dz9b0eTCXdsGgabGzK
loZQQplf57Sfra5eP6H8pvNZTsUek+V5G71bjY41PC8uBw8W1GeLG73WoMP9Vbk6qFLlbNVHGIUE
KI7+2hWyx6iLksMaJxxPui2QlAB7UHTzVglgw/h6U159VDboh1zjpN/2zbAkIXty8HjPxh/VhhGn
Ka0P/blTYfjb5Vbdgsh8Lt6r2INKXDN3XFMD7s7bsPjbi7q9s5CrA+OlOhRn/6GWCroJu2TaIqtX
PdNsEJpQxKFc9qjsVfekdKdw5Psi/cBLnWVCVKMkVQUz129z5U18Dwnx0ZpevWMRzHfDAyCtL5Dh
p1SgBwWmqI95IRGJrjjjZfKc8V9ffx3/+tASdFBVEiP97bZhFkCPqeQ5tGjLpWwtzTVoprz/JkTJ
fFuO31SdpmxRJig1aiLt478Z3mywgnjQrjoK2a4LAhF1bDJDWYVw4wPn8KqwTB1ytwHM1hHm9OJ+
lXP71EnyT5xAZjURfgMVGzaZJVhO/qTFZAIPYGtl/JBwUI5qF0y2QI13+w9kqz4Z59Q5OZgW/1/u
iIenc2jyAmj4FCcSazDR9CPKVaOPXVaxKz+Jg922CbApblwruBrs4LdAPvwCHaKUDiwDpiWtdJlN
Vc/bfEDcwOeebV4qjFJSRL75CICdWBU+ZX8eibrouMV1BtWOnr9eqM22kwYhxJele07Txaz+FxSl
GyTaDgiFFrQaM0WBAXyKT+q05z30yIkPHZlc4iVhq3YnBlaEjTN1nfqBcisoHnu6zJLbXWN3RIwk
Zfseu2ZMK2UYvLkI2k9Q1Sm69RfdRK4zwBJpuKRY698MBcD75E2zjc4108OtB9BE5AkxLzQ8+MUt
QDAJl9CmenKUpa/m3sIfAhucGLumbOQ0iJ/BhTRCRDTkqfjovlN5W06jZmWlQ88k2/0sdH97QZnb
UIaIXOtCYtFQDgrRieDAug3cMrk1AhryRZfC8+VlWuyWsI3z8OJQudSjI3Bj4eGVrwCcVPPODctV
QF3VvvSrWu3omTd+GGPXGSIjhdC1rO3S2ou5qDqpA7ODW3CEnW+PpB6gIoqmaDvD0JUg+qlSQdsi
xr1XmpnZ1OF79vCaIgbpIv21614saXqNQSbiDOs9M9Mp6sCn3YCHaXM/sc0yriDy4Dv8T6496tnQ
5nxKytSyTqA8I7s2Vu6f9L3igbkkLvzSBnm9q02Bx7lhtRZJjQo3MiNaziZ0ggb6BWvXiids1myR
0l8iDB2TnDjunqMkZ3aBqbXEPmYSWA/pGY6WtI1+vyaqSvVK8yx50eT/f0UKUXhMVOvaua+HZ8dw
Jho1NUzGcwAu/fusx413biOzb2t9NXBvbt5XtVvrU8qKUqF57/r2eys1Ua2fUvK7+ooMr8kaReOa
PgesrjO/HDtoGKXXaiQVrh8kFfu8WJjmPgZ6CPDVZUw5UNPouqpf+FEhKbw6hlDmqgRANxi2uSgp
kLCFgEeBRhRb9sDyLX9/ttD76y2jFcw/IgS9OYQb+o/EJfTqUKZH6Xqy8tmwkI6cOBJCb6hT5w2U
4WAtHQs1fDOy0FOND9snOMT8lIOLdofjlS7ZixKaG5J1br0nUAv5grAHw1zct2vi+rVxG27jS4qz
8zAU8TMOkiCc1Fe4DaTh/mdAZQLW74gGSF8dVzYl5iTvH9I4IwnPOEyfi4mFSlzvp6ut8t/W0wEE
QoIhLzj2CqRgAP8LtcRPyzd2hAofWo6qHa0D4UmcOrYaJSn4yNrV65oTpT7S/D29QrTz6PEDEtfd
ua4WmzVt5J0T2UaXqMrBKdBb3gWAiCki6d+NO/tjmRld6fPRcrVR6fXcDL5WtXvf/Pp/mcDFC6rK
T4si20YV6TSZQ0JCLDlZGPQLw0romaYnspWxg8H0M9AvmJW3N/BM+o1fHOwxtAWITwYMT+6PP51L
7Ia/dKZYwmTYxM7FtxwhyWVbUh6uquTHjfad2ox830Ze2djCLhIyOW7Qb4s5ZEOMLZfwUrKgXZNq
JOfnW4qV4qgjlY3ZnMB2G/jVlUIxPllUHpZtTYNTE3Kot/OYwzPC1/76HbWB8XkNdSMUICYbM+Us
zxn1r0R4TCx7IHOdBPywFHyLUB0c+t9UxHmwXBwBtI9LVAAHQFDDIuU0D8sBsnmzCGsabSAG/B5I
dsgZJgTiGjgfGjEyHEYI38CWxVcokHWTH07pz+P5y1vH+cKDQZPczkJV3reHis4iyqbZFaMbVj2d
7AjHCaBf0/hgZlF9lvpIqKsLQ0i5exAFuXY/gVINx0KnAE0oJRCZe7A7utX63v5KY3QWAOaTytBD
Qf0jmCBtJ4qdat/n+tcgDGNKGM0mowRXLOy7oPJrYeAB6kIwGEPlAco9SyfH+10rCnHAhKcEK64D
4U9Xk8wuinDOvfUeK3E4mz45s43kWX58Cx/R/KFz1jg7M0+OlzWRW7HNhdwbBMwk3J1/gvMoQAru
wnf1745KNtMZ2d5R3HB+t9kvL12dwKTiyYTRCikLMknNsRuEPkvS6CZZYAXYl8e1nnMs6zPgCCdD
xyl0q+N4VNCpNf9A4PomNW6tD0SGxju25Fh7afPxHGTxCutQH+skTvR66P8bCdRZOJwlje8KB/eX
RwaB0WNUK8Hc1cVbP30S82VvZhb1vbiZ7TlcGbm172I+YKHuYn7fSTU2Jju7v6j0xjDxMo2cdJZk
hr3DjxdNYJYd8OLDWV9ZDcw0Un9lfreCfezYbP0o2jZEqvWBJd10j9TP2UdcTMz6DD7qJ30kDHP7
8yFyyhBgAmTsAPQzXPZLMjMaHERReBcnqvZaCq40a17H0IJwv5vuXmqdusogozc+7H6T2RfYTbzA
mnwoSBRATH7/xnLtboNZa3/+qnVKa88MnNpql0fdXnVr+QyeaeUOz57raOcIcMuQN7uqGbb/BqQw
tVcKYOIq0f2CQ8NcUw2rqXhW0MkkCdqPU7n+AxiSduUvuUC2MY7TcxBlBEFz1LUCH+mQTb8NszLH
AXQEnwkiQJNNFpMTL/w9csau37LL4vIXcWOZq/KJsi79FlQcWoblQA8mdkmTYU1Q5hwJtQIc4GgH
MP7jHEFFWw4zu7WxlzUWhD8WLxSVkbG5QsJ0uvIEdw32544RUuvxEwRZxP5rr+58hKLAtsftzrLa
c+yetIM34CGsfZkt9QwtU1VN8gZzbH5rcfqLLV2CaSjqzuaS2TY4gVm2kRSo37PzQ/DnCCK0GJ0F
G1CXLdpFOvpucyZpl+YjHTmVMa2+uVrwbi/I38BeagYKwhuGUl2HsyyrVHikreHuqfpVSDWixr7U
MnAInYBL19h5DYzjlYqLQDS5jZXPXhuN7gLN70tdElRxTnD9ucfNGCOuFIQoYfwTfySD8nUbWaPB
43JnbOz9gOXhbZK2UlOXUMa8fdNYBZbQdeNmzzlWBc3fjBIVe6D77muUqKolTtCiRX21t6yjResS
UmPl94bOZoT160k71xF1IECfvgavsOlALNxKKu4Qbsc5D+v/dSkHWalC/MGlsvTRh+pxQE7FLntd
grFeckq6Jz/Bg8as8684lMrYkwqj9TGpwvt3zSMiFVV3ytQx58EJJFlfHAx87xawdr24HguRL+IN
Caa2Phalp8Q1COzckPPbHTVBO8NhgOW33UPpauwrkxHtVKnOCEo37vpt7YitQrEHa7K1bcLAlkJu
sphnpBEJ5YmKHHokYdXecUyklGzBa4dCT5TSlNWUWnhAjoYP7ZY8EUAjs1XdEbqArWgbZnyOF1xB
7xi7UUEvqzAkt7okatLjWy/bFZbdkCAkxkwOCvHZ/e0gkGNgutu84EL3uBA8fze/9I6RcUIsjqMQ
BJefcDDg5Dx81C1t3pUgMEzdAMGkv8XWlLLuHid+rhXhf/qgjFineCkmvBbJb3lSoV0r7A5MXORe
+KsAKUs1Pnao0NvY7hFmQspjwpUPNV9nb1WCjV6j1xFkDlR7C8ft7mLc7EOUbYrtL9tcFI+xM22+
hmtnD9gHg5k5o9H93rfhYDUj02TxhZOXUwx1egroCpqnJIeyhLNIdft7I6Lz9YNhxij4+t4CPXDW
5L0Jbn+mSNSQ8ru8Lye2UHsTIcAwiwVImXNVkLrwhtGX2U1Z4unzFBHBT1k+0jjkygczVoZXS0uo
QnL9yVWyQ9wCbIGeHgVLNU25K+Kdu8xioOnYcArd0YS4CCglozYToR2t8P94VuSgMG764n76AUBE
041Cs+DuIq2kZMpjPdNDCJKdU0YyN9RCv9aPWLyX63cQD8BHU0/pzrr9t4licQjGyWP3bdrrGbff
ime+oe47aK44zH4fqIss130BPeSesXZ3wan7YmQ37AwllrYocpJG2qPvJdgC3klB5bkEgMzSTkd1
joQ3esk13GPaiGt5COqLxN4bcxZjsK+KEGV23mi4nWS37qT662MfmoSQ8tWfR8K/CBCWOnnhNhOk
xIq9PAI0/FTNEXXEGEqx/Skt3LGW9X+cEC5dom5pUycUn0msVCvFSffvDrJc9rscExDin5m2pXv6
gc7iuQ7XvMFfrwwBIxxh0bXLbCm+nSK3u165VvbHqPwBIPN79uWIeRfoqqttoGSS1EKSqhlOXC0S
4LfGf2a6U8bTN50ZTlPbwzi/ZvsQMRfnMcQrI/JAhdLo7mAJ2KgxLeCb9CpOPIvAwztl5OrKRVSm
NyLWWPBsuJK1y8aAA00m7QbO3FNtIvBpOVRFD2ZP8GNB4XywuSPGwvZq1vJBkQCVYWrC6+Ss9q9F
3bLFYsIqGZOR4vJwSi2+tN+a+ZhogrrWwNi4QmaJrL3Y8cSi7Po9ILSMj1hWnZaqmRorlqioOvz7
JJz42/wq+3W0tN1SJ3iNFrS873IJZOg5j+017nZiUgGGoqDvUxkrPJKc7X5C6dVWuhZ3Nasw+U7D
A42sUlJuX6gZxe+Iga30AGibGjpXe+R5i/8u2kV5f7TPQcQN1PIR6z5s7WQrjhrcWsKO4JVmVy+k
Cah+r3gDqnvxKtfMF8xy7GlV2SCeo5DZPbcMTK8EAoynPIt9hx54U1nPTuH8h9F5SlWfgLlvXMcW
gPWFIrBowqss/a6HVo/wLdNSjPHwAVk5IL3ovm+qPo5joFpSR8Bpjm5FeCFwpHvnAtNL7/RIuVtx
S3r9+5lCy8xJHzxpIaf4T+a4DIFaCTGwiVTTrvwGBA6/8HM8Bra6Eo65YvDbhB7OMENzH+wGAvHQ
JyiBhYInwGCSqwdCqRxwQDLnCOqj9ks98WReT3pFP0doPzpwu4uRd5xsNs4Bka+eONqQrWTlZWxK
m4JBtqdGCZrqNAVGhNwe4O83/yxe4S0f0wi1qJyaWprhtUhivuxb6UGc9yHS02Z1C/ucWJMv3f/X
LDYaJtWuqBSiCR/O1nKH41BRboUr1qdEFT+ZBDiO0+obgKjJLGMEjhcfjm4n6qI2vdqaoLQ64kgW
vqgpJ1OUkHGpF/+BMWVqM1lXdN7x+PPEjeSdX733REiDzfWEz2GwIu7xK6SdwNpBRsDl94+SKJkG
MKIn1ZHrFA8xjk9MeH395/1SZ/+nwPAyBs1xVNfhT2UIN+a0jOy1obgIdHEpKlW6F7IBWQCjG3Oc
6NppgHcnrNqjJ6PeV8MtoPjTGWhFSdWBIGFPoNsQieRI7VLXV+5dzA1xc1OXcF+9mQ5tWNuUQE4Q
nV/IIHtKrQUyJqTSR5D/wnj08h9B5qovNS/jMUnsybk0u20KGe5wRRCwGNvul69g1w35dPYCO+D/
IiyQ+ufSFDx6hOYXD+bWItcGhbov9pcE0RO7gzCgHFN6nwuSYpPtFz0DiRwi19WvEcyG0NA7OppB
ABIZm3BmhJDgS1bFT+3bV5a/rnRHf0vF6TeaNzKbCWmvAQFx6Xgm/wNjZDdXrRtE1FfBrcCbXMu2
ogalSkpbicetCcZUBxhYVx5b9wwK10C+51EMAuSrwIaAyjU/8dPx53nqrzkxnofwqeoNt93J53SO
iLmVPP7O7dEfamTqkM/K9HbADNfeXbakYaCaS8c3OJxJxSLtmy1ntlX8TF3pCjBMmJ4hbXUvFU1r
2+VfHDtcdFBtDOFaM0WkcBVZt79rE3rOtu9A5EbnHZRXzGrs5HeHzBsxKNYYxRyOvg+3ZJEzWk1U
B+2WP1guMHS2s2JLMyOcxhNrdGfhcn6r2IlCROwdlv/F3FtRmFmNH6QF1M+l8wJhNrHhWQzgPjuz
cu4nSdg7L4GQ0WpN1C7ispW9T8ViJwiLbucH4+K9RLWLLYmuSw//dBC7/T8nJO8LZDGtGWC8CB3Y
L9lM+V6ZK47tfyn6tVodqiKeQoFaFZDaOf8tZO0hNzoYm9grtMSJcimo2okjRZvh6sirJmKLrGrq
mPPjsoWmhJZe5xisNfkFN3Awq7iyqwz0GKxs6Ig9hZOLdJiMKZEKB36L5ImnLaTcgPUmFNJKn0JV
m3TAY1zc071WaHn8sjr3VRMaU+qpwqZL7aGJJ09eNTa6nC5e7Z+VO/BzDuz02bNGLqsifrAQ0+0l
7Rulh3n3dIaHW2bNQEr5MrFXKxpviRgZyMKWFpNz81eE0+avxkGPL209JP4u0C6+PWfoDZj0Dc+P
OKYUEaQj/lIK/Nw76+QRuL+3OKik4SvTox4GyDUXUPfcWoWbNxFMuoJvd/U2ace3BI1R1FUEPs0G
1gcEgs6IHoeXXlJlvkqafGwuIPQWWEW71stRtCOgdeRcOdb7RVsHKcmfGL+T4ED1TF8HK71na0i1
hsAG2JrNoFLyvCZcizSGwn2C08hqpdIyZwORl4+EOndDFWY4js82vBe629LbCy5vrcCs1l31QeU4
du5XPzbt9HZl6rdRXRqjbouJa0FF4ogqELkoUtmF2tPiAxFI5dlxWBkQCt72PiSGWJ4DuHqTm3h+
pk1IPldrZXZjc2Hy1fnUz1ga6ZapOtbhsunx7/u/Sr1q7/ehgXh74lHDKvo/JZh2wgDtrBcxEudr
CuLpiKf+On7oj4MZQWtAroevvBP/na36jYz3HCohwBAc94BCqhb2JOyjG59qYfsr9mJMct5v5moi
vHqE0XCgtXcbWTMiGVR2mtH7e59xKQZRVHBleltrJtjZjUD0hk+li0lX7NoUqQD/+OywL04ZowuT
/gnlcqxMXTpX7hTSlODo3nis6lMBNltrPXJQyrtx01QSR1mDuEqV6Cl9u1aJxf03Ty9VxdxKGbEC
aVLd8+feNXHaZ+x7D3An5tA/uGPav1/9SzoxrGRvK5Tkn7IxKiopIA7yGx3+pLegouRc1syt4ESN
akwY9g0BqS45/RVo2gNWPn8Q/BI6b+l1gwqsnOKnfPEvvhC0nVkAmL6ShfSrJYuF6jSu6gd2vjQ0
0l/nlFdhXUAAI/ecKNQ5xAnvnNc+M/s7/XMq260uCD1daoGqupqOjHPfFm1jYLQDWhwujgd4C+83
1bf8YEzASPAC/t2a0aqE/v8DNsGXiVvISbhbXTDuwd3QEVp/O1ZEDQvWUZOY5VCpenq4K64hEHkP
V746UoH5FQ813xaZCOdTWDBi0f/w2jTMRiX5MKm240ILAvM3mGAppl1QCBdrQ3XRrY4Vp66hrbjW
K6D5/Ulnra6pvsf8FoNTXnbdiATBDz1IoyhzrGrNsH+yfVYO5IBYc+vynx0QQcwp4AALyHtsk66Y
+ThrAYsNri7X53fOd5CtKkQz118g9aA5QxdBG8aYvs3yQGEODSLtCVRcYWpYRauFVC+l4tU9j1aa
3Po23RzK6gt2a9ziJw1AMFaBF/EALNQ4Jyvyrkg00D01ovjhWs4GGAoNZtEvuUk2ZqQfPc8Hk7eN
DfAcNNAu7L3x9wJsVpTpzeez876rBTAI7+53rV/XP2fm1SkPoa+Yr+T8grAqMm8HmmanpaJz2sNG
8b9fKaLI7SRC2lmd3LC0oda5vverDERVI0reZ7hD1+kianB8ju6183fHXBqLjcjK3iu5r6s1SHDb
bmch+EnGzWD/OciWAIbZ4jPbcR/ADSBm+tSbUuY177KLOwFmTiRtTizgBS2CTy+0yq6+MddveXcW
23A2jwAACFt+XAAS+i5n0W2lSdjhixGdUJq6OijfHAd6DB7CrqI32ddsx4EY505jbD2osM+tnonU
84vK3N0C1hVu5XwbQ+gIWlgfUISfIDzFt9N+zym8OpFwFxQU30BZ2425G7PE3qTzYvoSZfGpUSST
+Z94gysVLC/7lTfwkOXB/9YgDYXdjq26u6XLAOqXmQS7HlAgW3B5fvoX0pI6DyFXmuRx7DL3tnGl
t9xMLqf+8jRAHRVo3KGjjMKGhHNjIyrNhmDZTBivVXVSOYw60pzXVp6OTD8WL2SDD16u+oPbl8kc
5YYyYpyqrFsiU/RsEEqrsLLP4ILXb3pecAa3Q6zjtdVR5skSp1kdMy7de109oNPhN5b8TUnQqMsa
iKQ+VZ2upRmJFO9sBw21AuhXV4I+kvrOAldJ2DeSZojXTVUUgWeQdjzYire8TxiFb//jm2JQJu4e
v0hpdD2ExzdGZVG6YLYK1cn2BH5vQxhRdg/G0agCx+P+ogmKaObZ64E+Wkzg/wo6oAQl56y5dMeI
oqQFunPEwfviyAUXy5IGmzf+0A4ocaRvw1Y2sl1NIfl0rBtnniR+Q2Htvi8MYh+9oRPOQ5D40LT+
XSrjwZ/rxEo3Tb8KD9/6Uvu2MkXGEN+vsRFtWhNo7H9p0UsWB13BbjcfcbXTm2XwVVpu5TrxnKnE
43dX62O/B816arBw9PD7q6UpoP/GGjtRAgDlegse1FrZBPutxmWUe2oDcO9RpmWFZqkpyfO48a3j
pm9V7CZ+J1cL0E60vtSK1JCr/2W1hKQlrV/QOyt9Twic7HSJZtjAQXlvaWJc9GwBK6eBC/aKhzSm
UcV964wGkJ3scICcbCczYosMznNGBoHN2BJ13bS7h1XZ0aT2eWlVGur5ELI2AHvf07butQ+yv3+U
HJvELQnrnXCiPTAV0a3XovO9Aj4gNEf0ya9ZowwvWsCZ+WmR+WZqht76jghtIQWJuG/viox7yDDE
4ukW4Z7PKKU5rcGIcfY8sTLtL6iQ0GPm90t61M/HHOCY20kjqn1qXVtwCECsUQ2wo8/7nDPIXJbe
E6vO7tOcKdDuujiqVyeNXv2q8XUOMVNR5cTMIlw+X7neySd7BzSbU2A9cGYYgEBjDg3oiamcUtU/
LVtArvYUIv5FGn3G9209EmG1VCLtp2s7JLM9OTLVuyOuYEFeDKhp64mFtOB8IDiGm6KhBBeC23Pq
bKWQUxTnNBBEFaM7U7uclIzICkZePXNhQ5So4MIVQf4YLeX863tCsBD5gFsqKQ69LMwC4NxUCTJ3
+AQkB81xuPtHjVoenoxciuZaEdbHziBrLTu76PLdMXIP/2cq99vXO6OV7DmXeW+nRZV2Kw55V/0w
rzGTrdIDC86SZNYziHlqypHEjNSPmC/a+JuVR/ovIPGXjZkbS5ci5Wa0LvKsFUGlIGdslgNMlFHD
A9bxFUmNQG71sR8ybIKv+ylPE7SziSs127XtqFKWYtFX5iqHWBGWPsPWv2dm47NSjsqoMe9bRFPe
XXvJSCmd4U02JLp14rtihdFMGPvLeyuotwlBWKFAGfZufnu5EpVDUUPcA8pr03O+jv5Hf/EsfZ1d
XZHAIz0dDb4Jov6XtmPstzUAGb7Tp6eSL12p85vCgSEN8ZYCM+krwarZKccP6GxiEoxdFowlIfvw
7ZmqxDd5EghHGZdqfTL77QuXPkXsXaK5v/VoTTi85QawWd5nnPiCd1wsyRfOUS5V8SUo+jcHPzoR
TyUYz95LNXA66OLQPgKjjxFLcS0vYGyAnArKPVjwjCE/j4B2dd/FN9O42NKabohN4gxYifPAVdPT
0O+W/OD0IREXNKpGz+5nwfHcigiScfJlkOgHcJ+6xCUKR2kjKFfwjVlFFPTs5eb9hawLHrKVDGb0
tEsDbixGkQvMyAcz/qdFn/RUubtPbx97dnusBUiv103FF10FcgsN3R+6E8DLAn6xoBCdjSaWYGms
qcHN9nP9Q0+KKCl1s946iiFfF2oyoo55jC/fMQVc3pdMQQoJqyNgL+9gTXu6AGpdBg014KiRSZFA
kQZrP8oyio+dXsGcOm3a5aYn+fWbm8P59G3uAVvQn0Y3HrUt/L9Yums4TrNisOvbuXfl+P2SFD+p
qRVBMd8uoj54TUgUtxJgz9ExTJtRasG2t8Nk7HsNluIbByjGRPJKeHwWYYUdE6AqyVB+Y+7N0biS
AbUM6nkYL9x88o8p+to5XUlOEjeXCdJmmjUYB0ge+xId95ir+WYe7nd9SgexcOkR58XjE1nG+qb0
R9GhTNXxPpeTRwqH53X5MdH2wBq54O9YAHM+u+CCv6REkapeuexO1380KOyllObUw6uXR8xTu5om
re92ON6zQ8OoODPoSFbuNaUpiZKvVrUh9TL++qclumCC+xDZ1zpdVSGiksGpk5gj3f03RE8u8teV
p43udLp5XkUMHDC02R0MbxOEOvB8QorR5Vlhzg1e5b+gavS4DBIyke3QPH7eBd8kJC3fXZ3+v7+z
eJhCkVUhYvY1Jiu4gHAPZRS8nOug0FYJScQFZbFVaUhjwDFsMi076H+ykVE41qriG/0HhF2OMrAo
YEyrNjLs42RR+EmqdjAUhKcVy/t2jTJp5WqHY/89olotpYK/Z1iM/MXX4fOrYs3RPn8zdWqDYiNr
FqF+Wm8ROtc1GlSmE2s7qTKDQ9lk8gJjzjkxmJxXt9afAgJM9dUrjxjDAIiOpyW8yhznhIixC37B
Fn8UfHumNN4aBqtp7pRUB0ZaMOERJu2hQBr8rvFTcHsoCuiue8eby+bWGjRhNnU+wRbZ5OEEIIeA
T3krU4cc+fG7+67rkQbjGPBnJT3K2REfLCFzDI4uvLd/30bSI4q92UNNBBvU8RrgvgU4kiXpUfnx
0x+vqZM8d5NWwlNmFlg3sAEbELbImIls9qc0BtBqLG4Vjpc8l5Vaty/+AwM6u6VGia8TyQY+W6wA
zenoD97k3eJtTbcw+grWZUicmZcAc46IaIKoADzx+UBvODfVzkxYsy8nrXHgRFCCT4hT+fDsplj2
4qpZm2bu+EutaHsw5sWF187LUEJV4QHmeMNoF06LQKlIvwRlZyWf8r1rIrbVNUgqx43qiIz937gl
+i4+pTg0aO7xnc1UUw9nGrf3T7PMUDM3GSh3RCCG9qYQph+nnlRUjjfc9CR2lHqMXGSVLTI6pf3u
n1jj7pYYOOY/DUEg1V0wL/TXvZ6as+Yx8TMXyJFsiFP6qIZ267GxwqQgFHmcV/KaBjWbVVrX5ZAS
mKHTWlrysWkli7TEiwttx1qXzHz/bRQmCCp3Vrluu7M4C6/fMoCCdq5E8n3mEOKRMv6reL1aB0cr
W0DLFvo8slaQUw0BlmKm/ZCz3f6eeXGLyGqFRw2RPoDfwGYEjiHBPe7J5dBn1n5uf5ixVkdz4fco
RAXgKswo/eoOY3ZGUjPDrRifEiNc5bhTaTrBzgVb5EiA2SMoMZHjMZThAtj2d8OhvOQcbAhhN1c2
6KxXmAMItuNjvLsp7CW3aRV6i+0Q7iGyuRNu+272voWq/gE5s9ikV1M+L1Gyh8YHGlgeZIeZtGN8
rtre5xgsd/l2c/Q8bzWkxRiO4wXPecJv84qRFsu029jE0941sCK1LrwpAXc2cROOZmC+bZBHlpqE
oIdUxAjP/4REo6G/DGz7fVdqVE+TKc4HDYWLu+zEKl3NeL8FZdrU0+kdEkr7WpmpNIXyOHGVODk8
G+OF5tY2BQVJw6t+m9uNN+KDUtt+qAAOHkuROOx8lr6Q9iHcaicLke0KW4RPmNuCLeZ32SxP52FX
3vMvD3lnCiJmsrbohwm5wa/rUuXZmNPc/SUV0m3KZ+4Q88z7YPrMNZQN2jrFRdKhGaM7qCzPh7vd
ve1N1lY6FLNpzvSDsbqigLS0V8qjFgKBONroWpY3ya1uv5sFVZXtoTiTLEu8Z06acZl918J6lAOV
47ApIEh0QyEXgy7OSahkL3T7b8vIwqxlGOdI1DwsBVxF/bNw8XTlXa3t6/wi8tPk2LfJ7w/z4xFK
fNW+7wKo6SCYgukRN5bz5U+9i9S5Shgc+sCFnGV5nZ1TCXDboLkuI/0ykAJwBU/aKz7KN0H/t+Py
t9OhDNbtWaAqQ8m0HPggmFRfPXm8/AAHFIIm2yctk7XMZwxvBC4e93DaXPP+E/r58VrUb3m12ZiH
70dz7Ho8/gDYjO6sZ1x+2JdtWiTOK5m9FMDz0fu+GkTQixEI6OlrlkFbloshG6AVdIuTsQzJjTSF
UnD1ncK/1jc9NlSmxRBdhGn8QwdLk4QJn+iwGGxnX30/TROBUWC9Lv0bGp2tAC6EBAxyQ3sLQas2
SQGvuS3TSL9UTWlrsspOxcxMLHoZo9hzKi4cXlWcT0hI2p6V7tlFDw/cM59Gn7KZ9kPmevk1OQtz
FQaUQW02j4McdG7zB2OsNTuvMDMI7d3xAfMoHZHm5g41uWZlLqHz/3S8nCVNEM9HuLC1r38FObiT
9w9CRPoF74YlEZ3//VSZgab+ODeVuOBDqf8HafnviJYCw+7TpGYxrDlJ8tvcwIRycMoh3iUNo3ot
0EjD0jZ75Qq5o7EeuYPpfvSDCgPBy79DtTl22NDxZFx2pzqRa5Dba5a15M/Sb/ZmoE7IXQ7Xqg5d
NkJF2wudUENGVJFe3pRbFpTFqOS+Lp0x6Rape9vtRLB+d0bjyY7FtIgX4iD2KdBbFiae1LOd7woc
Hvd1oPL1mQwa2szsCAPM4fRiYCHbNNXPjxVT4UlyEI0LqdgKg53i0Wz1pyYo0WAXzjfuLK6VaBb8
A1ezcdf1LH07EcsvR+YkuvysrscsGjl9ENBV5HWzZ+qZPDc5QM5/tJTJKJPedPDxJZxuAa2W0qIe
eVruU6e2QIqrxct8GFCjjMjRnxCSibPf1Oh4aNxKe4egsK8dfp0/GK6xfwn3C4bmQzo1KQJiyw1U
KNHiBHT9hYmRoBOG5lEcU1iGgQwpFO42p4cU7vIJq493gJBwbcSwFCUjnl3k4NC/8qJkxlw+fEa6
m0+bVURZDZjGKQddCGnjReK5hL5sENlE7S8eFhynpesEeUoUQz/PtawNoa6BRaNOfqjzltScfSrR
neK9DeFqS7dXmzOlHDzkn69Jr6KZsSpSRdeiTKoJmiWEsJ98uuR58/apd5lUUL95qqrQajTI3XYm
8PDPktJCEvEfwHiIymwv7ltiMSb+yoU3dtBFI5Zl05AjjQRj/erhRj6iZyQq0ER8N3F1hG+AkLBU
INhyuzsBaAW2qD3qa39JtThkUGeRFeFXBopt7qhZPJQN7WhfQkwy5JKyK0OAzZNm+PmmxMaFfQnE
ACR1xX+gMg6ie2QLDN/e/JAk1pH//22lcKxifduzRVGYxOIs0D4weO5lBo5dbM2q+5oYJjsv1ktW
DQsMXKlwMHLhnkfao5oK1c9Z5EjOMN1Q93/HoTWhucDDIkmLf8KOiyZhUpgFyE/TQp/xAlnoLhm/
vqK36v0amYogcazYyliMGdw1gNwcdvuLfv05wR+Zz/fFPcqw3WfyQEiNuM4q5tu3Aes/Ji9xkexE
+L/HvvWFbTosfWEQOJfFvoVzr4i4UoJYWxXDa1XmR+iBrWRHNiayosr0PMve80+n4b8uvgxLx3In
GL8AF/r1AzqZmaWvPEtVeM9efsBAkGUC4KOvAxAQFE0ea5iwc8fpxrpxbTUX6R0Xx22PdXB5ggdS
6ojHHGl8sth+a5XkfD39ZNBgmEFZMyZoBcLu7FSVXH2l9JBFWvkqAJId2RDBU/iCaOuhFErNJgQg
VVJqtWEjRKCQI4hDug/2p4Up+hLg5jyXoaLh1xjf8clKZAy0u8EaHWuVaatek6AH1QkrapYHwWwH
2vbTXxJr0dqM5+fuG12ZESdLkN6EKn4nqNS8O0TzHxoFmmpLgUuuA3pvXm7UMW7dSxk21XtzVCrN
/8gydmPYdYEU0OREMiazaaIazV8W/l8Y12U5S6zZKJ4tj2CGFfZLdPRC5AghjWoLJx0jtNM5Rns3
ZmEMfH1nERNXqxEyTU2sIKpbb97Ly2mBpyFir66TJA70mi25P4hubM3wcqamABxRgpj4PDwSu1rg
7LDdb4LguBy77ZN9DsBo+60aN7cLwLlC27vzwpJ5JpW8vGc/Hif9b6iqNhOh+698wFswelE5taSH
gEJnQCk1UNbZ7CUQU7n2LDMIeoGPVdLJmEJ7UnwQnCbx8XRGWME2dHO2HrpEuokTxeg9By7DID95
c/rx+wEgslOkVB6ohU/CPXotjv524rNyKy42jzVQm1VyQH2ZXA0GcUmiVPlJrFFbrL9e3kA0b06r
/uR8s5QY0QMJkfxaJnIoVILMlqx5dxU5k6Y5fxyaYG5RiJZEBBBxQX1ZuxUgUQ3nqs9ocoJzVCxh
Lc6U6TR/YqB8pQ/gdXFT1bVmPcRfwCirw9etvuHV3ek5loMbUa/S7WbQK81dZDQTt28my2ubO1V5
ftkZlyzMqZlhWSY/evTtYloYm8m/phIvvlqDw5dNNY13EE1Xzv7bRafDqeDmrLdF9d/Z79j9r4q2
sllsWFWaaw0tflx9SieiJY3VfkP59K1OF7QwnSj3yfJhb50366FOwmSzInf2ld8FG2OvijNTE5ZW
FmXYxgieF6zbDrk1oD8xQyB6L2WuvJ9tFjcpkizu8DFNvHtrVq8YgVE/usk5DfM+zS7uM4iIUm/0
Mccy415kEvXzyYTFPLrJrqFA1pvw3bXxJoVhPl/wCpiv6066o+u4Miy2x5BPyeKR/AgskCkLwAeK
9CEm9GyVLC94BPI+D6tC08g2c4h9mzB+rTF3xT3y4G7t1hkiaSk9MNLqJCnA2BM6rK99w5WE7iTi
eplnd6A1ornNWnMR09JuBzcQhNX3qFOJbYioqZ0ABX9vjoFhKYcqKE5NxxMr2m0uXjCdd+TXUY9N
lr56dNBymxAhSkblAh2pcsJQWivfuIRzwQJp3K3RQbShiq73BimYz4evau1+rIu02eRvDu8c6gKs
aIgNaEkF6f/mywObbIrp+klZaUJxITsXJLwBTXyyfxFh9vZHmi42yBfc3R1nRf2NgdUR6Fi90GjI
hHNjqwH+oKebskijL7mc9Erkv+9m6p7avcdRh0jr8Y4G1vId5k7N7y+BKXYph/F6sATHEJEsXKNm
/QnpsGFKdUp6v26rytkqQs4mH8YQ+AhZY8GgD0rpRCyddjnfUpBpHYvBp3an0rayEI64qZ4RdA6e
sadoaRDg+vR4AAk1HLl6nNy4P8ByEeiw/0x7KEKsU4NWL5yLAle8Ulx+6NuQat7Bo5Lu7H9J6fS/
nQFbwpyHWGvFq9+SIvQG98q6Z+Ll1yv8OejUeWL3kaoxTlVKNaOqLurgK9IAUpPEfVFpNV9M5UIh
t3IhvkydMz52sNFQWfsHHUDQN9FOsaUMAgRT5c3fyaoDBrCNxH58XuQxx6AA+VOqSGe9vec4jaPa
I+GyLEX4UPBiOA3HXrrZ/zQpGeuNOmaVGJAEsow1A3+GSii0yv/mWQrGLomc66U1RNObarFhsu/7
ZDkaZqRtvIU7uP3ba2NfCnsnWWeP49pJrp09Qjl/06BdjxRxTRJj64+6mGpXL7w+DC1M8FwPXHnn
4/nP+2sb7tMDkRWsI1I7hnUn8pPGv/CLcvACHaT3iifi6rfuHdbTTYoEm09Zx3puqfBdTt3fmVW4
Mr7UoQi29hPqbtFTCRE9sOlkdxuWmrK0LJYlasOVzvCniblFuUEjfNwBi4rRCqVJSDNslceGXaxR
EWwDf68AUPhM1677xeXfhuVhMn9ycVgYlOhGpgMyFn0pJY0hTOn/iqE7xVsgwiY+WaNVVWB1RDRO
95gJ0Kt546sFbm2QrosWOJl8eIqT/G/y4IL7MzmhxqLgHvqtxEpz0CKON28x1YNk9HYPY19IlKYq
x44I/9d/U1GdW4xDgyIXi3tx5HrcMs0EvFfCKYHJbHsuL6VYvk+TYxj4L/De34yxskD+MBpNNYX7
aVOdu5Fc1v1yXumupehX6GxdnEEU/68jJ02E5Gge4+rQZH35/Yp16UD1jynmT2JjCJD4jbsrvG6v
ehWQTWNuWZ1GLGzwoqKlieZcMli3KnTZ21aVA9Vsa/X3tz6Xqu2aLzJd0HYw63GNro7HuNZm4YYs
NH2eu2H/C2TodfF8nDBmJ/+y2m8MfVE6Np70EGMpNlASVrNMCpEpS4M4aGacaLWz8ny5Bfe+zSjZ
8I25c0ID9RKEniinNbxfEKhrWV1PPOQVEP+Fb8kpuHQ2Y6tjD5HbgDDK6ArC5HV3eswYoV51zliN
9qRcPuYpit0MOJuFTESp0lE3pzqATpLiF/Ph1UwB9e8RHom6msrFLaUxBbxUPHphsQ1p6VE5nhDr
bzqf57BI3rTFuPOLaVkD5s4hUf2J4GmM9DSHgLnSYj7kKUPv34bu7FE4rXvRRX1BUEeqd4FBrbmD
rm6h0hP25vWtEFPNQD8Nde0Ob4ryFMxnGWotuQPxGrPNvCxKpMs3/R503B14gxpjlAEcbGzcpgg4
AlVMplHlU/SrOz4SDBdn/py8u4hx6IXiuoZl/hGSc/2BqVfj5/AvkUXEtr3MWsxljkOh136THdm3
U75TuEeqXhi7c0Lx6D6QEWMV7+3FvVKJ58SWfUJvqjl/EE6Zg+u6HQt3aimK6/J4sww5wmdzCbQW
qca2bvWWj8be4FR0upyQ2Iu+uY7pGAhC0uN067sbDRmoqCRDPtXXjeGAh3hJGgt6w8bdo6DfUOqd
tY7F2I8+SxTXLCg4TRgIcXUod12X8YPjiHcn9F1d/kL8daFwVsugJYEpKWOscGG9RArLqhPs6544
Z024eE1/WsUTqHcvI1cliPVwhv5kDypTPN740DL0Xr5TfQXJF2uuZ4uFTVsaIgp7hzDlM1Jj5sT1
t6lWxd7rVXtS8c/wD97gIvUoNjzpYx3jJsbVmG8l5hrSoqNNtMqce3t8hEwNt1nnS46N0mWbvC6u
3R2/gl+4/PqUs8r1JR68GofhGHdk7eM5iZq/r7EUC5h9n3sKcorjIYGOhSlNxFX9ESEwaTJ8ThWb
285w7+3CxCrxnkYYpqK7aZS+nbGKvqPNpB3chO3TtEIqQvYPDyzrnXdGrGKIdIqhgzjwtTlbwlNH
ysBYJ7ciuoMMXTzRYAs/1nRjex0DU94i6plyw3YCsQOYrEIhpU76IByr9uwQHaOAoyoDp1p7dxH5
+gz/DJd5ZqXxgkjV2xLl+xgUAzbsiamYNxzt7DDqT9ozZ6/fTVvwqIBvw5DGibp4lWBA5C3oLCC/
EO4r2aYukmU2PiU5xE0rttAfz6vDhuvFRoPRB39vAcCzCD6rLBJxwEzh1cY7ZaeMHf7sg1rI2STZ
vdv7VyDqeyewEoz0HJ0K0NSpyXTF6k54tktZ/rgqb+jIncN2EGJSy4DhjU+Y3qTWB3myD578VhEO
+psSUUvpv2XBKeMbaJG+1lsyCF6+6jJjzHJpLy27y01SAXnA1V/jIqIZcsZZCX8SXprxEJAI0OCm
xPw6u1HV77KAsjPoH+9ceSc5evRdDctn9xwqlJe0d41QSvkcYOipT7FWmt/0dlq/2HmfPXF4B0H7
4VgW1qaCdMwC0gjoqfFJdCeRy4yyRLVR/mXJUZkYSlKvOJArxJ3mehakx4yiMLABq2Pt2PKbs7oe
tyAT95n92eRAJQ7IVG4CVOIvyK4H8uw3P1RKr2zEkQ2Ls2XqwHiavRdD+Kcu9ILRCafygaU/hoU6
lQXkXDVA5foSv2yoYwGFM46Y/YKujhEce6KSViElPi0xeDNrR/0/1UvzqbsCvhSXJrQvniKhvD63
3mQyV0UKVmOMeWD1GZa2PEIQMDq1IlZJOzkgfOQ4m5Zwm0m42kqXafyUA6Kd2pp3FmaO0BjNndSa
4smXPaBKax7hPyJDfFVpYRIzwP8Y2hqHUhD112j5ZSYdEc13pLCdoxkMPCADcQ4pjsXk7/xHP0p7
G6yHvKeBZt/tBYkJWEGhxuPF3Neuha7BhI6fRRrPLRifPCAJGm1WYiGmjp5zIYF5PCV01Er5+pEe
QhpQvvEKtnj0bggF66MmFep6O1c/5n2md8lglXbwmPDaGqmMWfrzShdRMQOvvYuSOPmxE4CQBZ3v
Wq6IBZFqhs+cohNzNVnFObv52wL3CfJ80dLw9iKa9ImXN07wec7p/wnyaHx8ZFBwEMXTuoV9cmxG
P1cYGMvis5krbjae30jGmKWidoOgtsNC0ClGnkSU9+Ng6eO/WrcrvaXuBOPaD0Or3AJhu+Hq5KXE
3lLuUhz9qLTdNVDlxHVjNXvQa/NTGSLknKQGY5V7+58N8gWNLhu73LP34wQB4PyWTwt9pHr0cy27
zORlxxicC/HfnyG9mXWAMyttZLlCAkqLSSusogGv4/SYbAv7dU2RzECpcGXcX5dGIBI7BmAO02Ku
fKPX75XP72W82ec6J+CdUticQePChdgGA8E5aF32dYY3EPhyDUoz/2dBSczDLKWQ502GqaVKh96m
sqKhEda3JIjAIxMX9c8SagmuUPneASs2Zwi45vfyJoqVSo4sbGbyV+3aYvWsfk6jwCyiEIrnsNB1
S6btmqi8Un1TRfvCbl1gDMpaGeU878n0vE4zz2NBevjDGdnNBSKDPlJoTBagjn0zabsSStZjvgub
oxYqDyRRX59vnAVL96yoSYdiluvNXnFpaTxPazrOoQYwXgbonE0HPbLItdtLXVSlJcTI1B/aVaKX
6EToX1ruv7CraRUbnsMXnsaNMVMRk3tPa9bGVIiuoKvUdYlwxm2hAFUB8bSQjvX+07s5r7hFOOab
AgXE4lZ3fkzwT7DycVEYqmv07sIyBvjnmgHL1Jgav7mG08r9i+9PrVLKnMilHyQaLFn0maVrOi/W
2OeGJSwBE/kSJXmTPpBlFFoTyE1BWG/zZikpn7HPkg0t0HY5ixMjDhk8ZF92ENxrB5HMm/IIl26X
aoU7BxpocTDWtmt5oJwZg81f8+GO0v58HgMKsAj19L0Syplhx5Qb+aABcQ9gfI1WylcmKF1JBHwH
QQyQPK5PZXaZZH1njLrX4qZadahQN1UyrIvmDWzJC36NB2aKUJq2Z+PSPyAIRln3OkLH8wuZX85m
VD+3G8yg7Ssjm9eeV6XGJuJWDIEZJ6UdQKpfJO15BLZ/HBUZEip4rKm0sNBkJhW/Ty+Ybyn1xY2E
5RYwSSXtarSsXfdgJSflfW4MeonOMm/sMCC4RihGOnimHPII9XcPKt3OSpRGEOcTjvzLXzlG712M
dy/JaU30AxPZyIZEKKSJ7ti22LpzVijZfBJhHRiqqWZDH+pTgLi9/6eG1OFD8Jd150mQiI0FnPJe
dSLqQYzCZOPS8ItldfOhcUQAumjqgHQ4K3K8ZXvhJ5AsAQotBAzY61DGlUQYKSoRQpIuaQxWJWoe
XCJyLRMBVKoOZwujNXrx6huLiSPxOJ+E10rJKVIJXOwgud2xqj0xOXg2S58/hOAnuRQsz1MSqqVA
A8ZQl8ALGYv8aO1BYiq1KcmFT/RYpOQnSbPhYvLZ/6xcOm+DRvzxcUvLklIdIxZUbeSZ+9Z7n1Yv
02Zb+GFxgqyM6S+d9MKZjtsLcTKcrnWpbyuWV48c0VpGTWMhGnToe3ug2d7At0H1ihpHIXLyPVgy
9MpYaO+YA/CCP0T6zGWg+hqEsWsnc9CT5OTkwoFVgzSe59w4IqCdhhguCFy60oL1PCMg2ZIDNDdl
EBA8c8H7FhAkGUsshP2/JkdCOnp+SMZbbRzpvVwz3NKHzFexrwwZ+Dc6J6drldUqSoZ6HHaj2C3R
uqedACE0L7vjKTT66ZsZl5MFp3fVaVDi8/9pFAjzvBU/V7VJZ/rvbwaeEDGvgtwa6qd+v8fgr6Nk
BEt3o7lt8N1WbHQnN/5RFN03kFhnB3hdiYfa30WuCUqJS7wcqvbky10iymXZQ0aIlL3fUhUchUkD
1JaNbU+q8vYrSEBJk9d28ccip/IPKg20j9gP5c21GA35RREO0rFZ9+1DOC8mn+Q371djJFLgHbEK
J7tTo1OsT7+9S3nt6lhPHbxUrpOpIB5JPhI7s5ajyX/uLBN8ocTcssmVShYMRAK+5pySXu0RpimV
BTo3xwRlHfET7MEpyszKwMGGPhWtohrdRlBztyTbrvbgWhgAxrQ+SqnfIGvhKtNSbxSbru4Iau3W
bVxUywJ46fthowFo/q4hxD2sYwTL5VHC3cmwzJ6A3Z5HJcCKFtGzZZJ6ccKac93moV5GZxQ2ehyh
/mj3VaB8Gd7Rr0XoU2X3P9Sv5Slu84+rI6z/zMAHT2djbtrFNWK5F+UBh8Z3Wpj6xsT6N7Qrx96Q
e7xsDfR6cvVKZYmqWSYvjVrQd44g605M/yHnzHKyYQqkjY5DOFi3TMMlQ7OgWYRCqCAFyO5VNFPJ
sYw5a0FW0d3Ai1ynmvzFEyKbWqT1tbjpgE660qOoAlXh7XGk5o2Sl/WEiES+fz2NICk+oFppHSF2
x2ErqtI9M9dJDK3TVPng0tYgXLcRsB3DTO65cm1Ilz1dg1OAkjAWjlFHRPwekqGTy6VSmS9aMmG9
ZVZbm1jlXz83jQeek2Zq4wv0/OIy0bn9FHdEjd8jSAFBq9M5f37DMFpKN5BSGwf92hF1oCL6mzYK
emqsQXCGOCjYRMNE0cgpTIC/aOJ5f8ramAHAv8AkrxJNNJYMOGWi0VZZRc6iV+j8qwhmwHiDR0w2
5w4rFHqlAWOQ5T6EemUnIlDtHkwthzQarKI05Zta1jjNA5H2DIV40VQgsfWnz5OkolWqigfJHl+Z
9RRTj3lQ4lSWhAs4rAZvUBf9sY8VnfankBkgThhb6hs91yIVvG2nZpnI8avEyBymUK0Q8I72lo2O
tTFLi/ogzDNrVBCDthNBH5XVsV9gw4x9NfEhLmn64gYLalWWE6KatfsbpZT5sdxfdZqEX7ozCfGY
giQmAONNLvsCmmTYLtYhLdmzJWS8q+dFDfuNmlOmFSmRiZVci7hMmEYZ06Blagaj1Bm9ao374v/q
BAgBsofxsyKBgzXdCDHmmuyBx4lgEoPY2N4Ekqo5gwksWk527tlqJCnW8wrTuAB9obSpwNe6fLKS
f99yDqTKQtlElEqUgyFXfZ9mIYDxLA+JWiPC+HkA0GkNgjSvJLTh2mPEpLVze5EunLQZ8xYZ/var
ospvr2oTWrBeqQxNcBfz0EJgWldPMHg2sdzTpTvY/Mg59dMtY3Nx5KQfT06uY41qKM1HXUKBkB58
aUc2fY7mZKl1Lyy+GjapH4FbhX3DSTRFpJUWjZ8uTmavib419UdgKSG6PLEGVZEnOULq+uFAB9QJ
x1n1LE8Ac6PNwJ/+IhNsIx/Jgbm0HV39LrdoUU1slOnbo0wu2w0L+PTwnp+/2epOJabVeYs6ipy9
gJssmd4E+qwdPOJTpeCy7dylssf44EkVirTAybfH4kRUY3Bbh2QojB2KeGWTCCJoxVguNGuRC9m3
hn76wr4Uap6mLrRRGEHdAu34jpxyxuPVQ1BdX8l+mLzMdLRTb2r687xjkeNq76IqF1B7cCtOdmoe
FAgf4g4+Fv7Wrso+ZifVdfmuU8hSeEyL7BybAmidh1/xjf2fDwCB3suOmz7Ikx2A9B++Ulwwipfp
tpoRVY44Q5GGrEGslcnraYv4FqYTGQ/PCZ+ULhFRTt7G7h6Pb8TRZXVKsT3K1a4LQTSceatkWxsp
SnAdhl0ed1fhrNmryJJwuafcDbgLPvtLtutwmRFgj6g9LzrWOuyZe5UB1fbmdoOlmyHhSznbD2vx
MKnFZCp1PTvzIKl4lbEnoyMZ4iLIbkN9ZYrTcDCmIYpQRqX4KKDa5cFdGX15RNOUVRTmKBfcmnmU
zmzcUWkIkM7zhKw1PcGKxT7SYeaX+YxT8MHqj5rQmAUqNvOjp/yoWPQwIUkfsG9m8YVJecuoWG93
FCARI32U58a0qvDZFCQMhINtKY5dYFt1WUM1VoVo/cWrumWNwG1t9+aZvisgq6gSZJvyuvkzBGhn
0jtQHS7wjv1FEah84lDMSYm9gT+2gOAlP5okFkpqRLXe1jQzPmzdCO/1ZdZ7+rGHHzjSnhWx/ODa
AixCvf1JiZMRmh25M+WDzl7aYAxo3OO+BB7WmESFd/tUsqg9e9bqcXTJovK/5psil3uHpInlXlmB
vn8VBcvtjTUW2lsSgkLm5E6vBrSNjJBY60rS6HbEbskxuniKbOTFcuRBrhTXVLtSxAJ2/FV36Aum
8wejwykvzpUm4UZbgY/qhQnJTybnDrEx/f9944yJQpNZL6d7rhDtRrtNj1H0V1MNfiEGPmqM5vAo
ALxNWo4V5AoBZzrhejQPWfymUCYPJd3q4alvwBeoUaOaHBK4DMjOKkNy0HGY4kYInH0ZOo2f0d1A
tA7ufdUwyqrfRwb/uBV9ciIN06TRZtbId65taTbsoJNfpUuQwMyVNH1U1svbrRlE13bf0RchhU6x
zFU+cvQWSTidHRs3lXqNkxdiKKdMIpAAYrZf2reU7FSe/I8xsqV8kLOm+1VYWES4X78WhLCoBO01
VurDpFrc4+fXThwiQbYPddlwkvT3+S/i8cn/msubmDPlSoYbncWBHrXU6US5ajl4a+3rQq0kmGOh
OquFI7BtbtwcDiEjxp6y5mz8LAA/BKudw695psU6LCLV2msbcgxjTLC07BeB8/UH/Jv5Wig+GLou
k69vMZLaC0ZMU1rh9WXhJba0aNLGFIdHaVUHww1WvCto1zivh1m4yK6ewASoh4zVK9XU74ieD2e/
lslJvroSPmm3M6e72cKkwjsYaaI2FVOq8OSDtKY82GEv1yjdgp6LL2S5jjfVuwhNicbL4Fh5gNh2
LQX406JMPFjIHS87gm+b1kxrfYOMr2cdw2oBs02naSyJ3P9mhe2FTIABkf0/S8STwEDmOFpTXQ02
dsrsdNAqwkrbhilRxtMojrs1GASN7m1xXBt9DWGvQVqN/ml16VLhAN4Bp9C/iaEgG8Sn0lTMCRqJ
VRWLJo8+hj2sbEho1xr10Yz1Kxu/9uhhBn1n5GNCEbWzNK4T9XLEGzcOBISLiiqM/QKfRYAwN2ep
XtavCN0C9MIFWNLEZSUWxeQ8uJrm9BaEqBzd5hYMVfgFp7H6svVeQATOK5Byx7Sh3/eKCV2PQt+6
mPbmhH4PAThqhtJsN458vmOGizS5LsO9YqXDSUeXyh8LrZ1Cm97BMY4InIc3XPvGtyZAYpU6/XMB
4pTnPysJa5eZdg6MtidOQZZBkLQsiEIxYsuoadVhhZs990u03Wb5cDFjQHi7SVaJL6iqTDyVd1G6
nPRxioBB4JTd8aS9Z4mm/NZCAW9Kbe68GBckwRVxR5Z24lD8Nv5FcoF5PU+NYvFNLqL9gZ8wq3xZ
3bKwu9wSpxiNJEZtSHws1hOXzoj7rbXyZ+7bIMD6nFT9dmOBJu2vYjFtdVEHFMn92xXhiQ6AcAmj
E5d9xU7L9tUgRy6ddjt3rX9EiKAYtXiM5bh4y9pv3/kn+F++2Tur3/R8nu8aK/02FGy0teqcFzM0
ieN6kvnxReHLsXV85nC83jmRSh38MOJG5h541QnxN0SX370oHJslaaR8ZzWo+q9d6nm4TYMlYJrR
xHdnmgNP9hlmSXMO6XdS/ahdX8qMyIFhA3UBJgTDT3cWEUe/UDzHh5zne1D7LNw7PRY6Hn16Shjz
cGUlCBWldi+ozF9Rto5yVmKdjQZqL9riBcdpXqWPLn1C6Y8E0B6uHIIxwI2E8o+ywelG2MBNfACY
R5ooUrxY+ByFhUkJqnvvlsL/zyE7kDbHkmHTWUZKVTWqJuRWO1HV0v3XN/8jxuppdhVQI5B/DS/y
gvWEZ/zXX5xfmovs/LJFDQU+n7jaISEeWrua53aH5HQFfAtA4d+3Wg9PTcR70jy7WWNNhTqPNITr
7dX8wf/aXUp0E52s9GSFfMd9v+2AM9eYBCMuf0jTMd7KqyegwjFb10j4PcRotfd3ElGImZXuZ7iZ
bOAZ+bz7TUy3PrMoFoV71pA7p7bJCy1XKojvY6Vu0bb0J++BqiaeewJkbEdaqQsvwy6PNkb12nB6
Le+EFVmVQ7ohWlR/jx2A8sZwOc5yDNVxE5CX7XfMF20+3M026Y8WArQ8niN0u0l+t/gsCXCtDHob
DQ0+4Y8pv7r8C9y9UGdzDveGJV7Nprn1B9/rJdAzn9FaugdJXCIrpfSTjfSIzXfQ8U00Gc9sHtPV
8LiZnuwcCoCn4qjUW7uQSFl6m9fXPnvhJg46OE0HFFMkmHZB7TvGbFpekO3GaJQNf47A7BsE/cnd
833d0yD+RBpjniZAd66GrkxVu8LbtIV4RKkNWgPGSMIr3AbTFW1Zc39qqpBXCleP1qsliM5IEDW8
q7cmQp6LofOUMlBSzlKRQEFRLqDgyLQUq3ziGFNNri1ZPx26zWt+TFg2daVOwCJv9dGShi0ILJif
FNKkxa0q+G8+4CY4FnQWS6edlb1aflimaWhbHzBk8P1+XhBaR4fgG1+dFpAuXb70ukISE1bVAYD6
dqLGGFZEa0k7AuKpAv0lcwpGrGyPsCKzN9TXDFL1RzuqAm+fJrugOwj7MMhCFFDhO1hhxB658RS1
WeP9raJWzB7BNdXF8L2bXL3kRn6nbAB7iGEI0sPSoDftOkambTVmw3uQu6un8mnZK0CeuG0LxOZ0
oDdTFEtqUxOKBbeLpbt14pW5AuDkdoD/4YADntmqC9E88nfFkakairDkCp34d+o8h/s2i4dAfMHn
VGnhet1YW36MDcLYEtLup2AsiVON8tJK7k92Q3i+DNWtlYpp5d451GMHfdCxJY5SpipNoensdr8A
46aVP7I6SOjZFLCauz2vFau/zuzRnYcB1e+STYx8wjFLyp7nbKp+EgmS3WZ6090g5gX/cpPrAeFn
djZU7uL8TVvuC2ImeJwZm6XDIBvAuYsl4/egCQEk2pPiI1ipQPA/sdmCLnafolKb+a+NIYCjqbFG
D9jRByG1ZbNjoxHEwYD7p+BStL+o2Vlw7ru0WNApoUnbOXP/2l4Wp0xKqDAChH7JK012z2XoafUZ
Nff5xnvzW0ArMLWLxMDhczd9ZiNAXrFxgPUES+2t8J1WwR0zpgBGf6QiAeTzJykJSJ3db/KqytBw
fVAviSUeBJHqViLwZ1WodpL+dPLjgQ0QPaqq+vnfyV1zil3nMhujng2Q/IhVHtMQBJGxjqQWmj0E
ai1yoxBzMpcvFkeMPrSGv9GyyI0ka5ovoBkWzSdd2mHJBjZLllA9vkQdxs4QLmvfKNUUJDrSqZtH
8PpzbWZtMSAO4CZVm35LRKTVdmUICWLNN9ziXa9sVjdSWr6RCCl917illpvcm20xavxqRpKF0Qex
zLotZT+g9yu6o/S6hDCg+I+iutp3hlSp475xpx3jmqRmq8LUOKm8HQR5C0Kxi4VPW5A+BDNr3tNu
8U7roWrC+e2T5NXjh41m3d9t37S85Y6PE3baD1nqJ1L3mIzcXv13ZK67DfYzxKpbuC3SGT6BtVQW
7RKCqtTBBU7aGOk4ZHx+hy4fYDAV+7RN9eAswXGoDgD8d03e9x6XeUoul0pkJrqnRP6REdv1jIWy
eVzqObuNB01BGqilnD3JUaw2TBpOLzT9AykRFA6vxt66qQOMXV+n0vxB983d556vuaAJxYdAGM/F
uVPLQT/6NVCsbnEp5z+BS4jpy2zY17J9Cxf3oyfTyosGcARYJrilHh90eS33YLEcS2W8n45AvFBo
ReKvtzedzZjmoK5xDNAZ98YrEdXLKiT7A3aBsjgAI9RIQiSz2FsCgWDFlaRGGOBdohzyRgAuxT/L
npG3pBGzjTY+O0+ivp0GJKxtZ8obCjON7fmYt4dJ12U7ZHRArgqaMLpGN3JJFPV8kSisEdpOelQM
+LF4M1PNqmGEbNzOAxCtN2r+UIjffNlpiYMha82yIL8rSoSYFGovRiodaQDVg+u7NVuELd+IE/2Z
X7Ei5ZzYwwU7+d8sLWGhGsLZSbY0kQpbXJYgtQUgTQ3+zEy+nfuf9i2M/6Peg6MpYjpmQefS37bA
mHzpZWRAl23F1uhl7pumSd+7QUOPWx/2y90ZERuvO/qhOvieOsTtzYA2Tt82M2ar0oX+VuW5EexF
3iRvrawcT2yZqffjCTvbDjMNt0cueG2KDoIGe4hd4W6KDzp+2xrERqF9kahHYhMDblL8Fzmqp+X1
kYZYV7XYLg7SsrFFQhqpbQw/1eJm7lL6fPYaPAFMVXTBNJ1bR7ASQmULAgyin7pLQ8uhCswOtpEr
tfU+DoXk4PyYz474kQt4uAXaz+yWKiUYnqIbFqH1VMfQThCBxzfNYJEw9oP1iMc1fCxR/ySlqs+h
yHjBcHMCn9T32RorkLn+dVc/AD7OZ+vNrBfea20acGdzeLe7xKPK8YS8qIBPsUNTGRs2yQl0ZWI5
lM9WJo/dKHxdZvKfuQbydc2kQqTnKk0PnKG6A7ixVnYxit/G1HrPAmRCkFeINTVmllfesj5QsSQK
I0qh8U1HMBjSAA5Ra6/T2/2Ppc6T2CKt7xHLhnW+TBFr/LgD5r7/BIHlBaSVH1iKRAmc+Kk0XVxc
HTkSs2NvWpLyO0wYtpOZq+SpOUos35Ktb65t8fmNvZClkzVyEkqGES+PM2H9qWsoOJK3NW45G4EY
rmgijtw6QYO2UHa5s/CIr5EmTorSME2ajuayOe0D2N6UOIYW7uGC8bxgLUTubiGwExQLx9SI/wV5
+rJZ6TeTtYoo1EA0raj+UVLDXfWsdaHc6n1YL92iFT+tPcZ7KE3RdV535IaexpTqnP0RiWCsDm+P
JNJ0izwyRKwto4rTYj1U4NQJDgOXRIN32Zuccgcc1gLmKxUhq5gP9eji1BSKviU2t+HDQYTt2r2X
iTt62xY4LXOQYGYHgB3G7FLA1OFhPbSKaToGcSlVsPS0YkZuZBEQ2uO3Xe6bWcRKUx1yxY/v2wCT
/coCinh/XvFB07EbcHS3FRThCkG65J5Ys/+CNGcGHk3Jx3FOOOlhgZvGKNBRD0XFY/e3m2VyvLkQ
JAZrdW1J9MgrpLsNUU7tm8B/a0Gc1S0rrWDfyjVc1ErBXTYcs1Ovy+ErMKnU58FjVeSUqcrSIjXW
Af2xkCTrVZp/WbVGIvrx5g9klZ5TyTqpMWgRFBA7QFGDHD/yPlYBDYNc+p2SoeW891bqdNk/GuqT
fwbr6kq3k3gOo9SlLau3wprE/IUS+fBrt4V6X3lgSqfVQXQVbaP2xwLEQYWyioGNE3St5IcVdLMM
WLKcmvZmJXmBQP4pYa0w3EWiaL2GuDOdXtmc7NmXFbrBfYJsaBHKduWTdPik5awK1XoId3bhnD/T
adubRubf91RE73qyQwGA1OkFgLRwAYUhKIejRTPXBtY2QCYivCGHwaxswyBPe7cDUb3vdskUmans
RpAIqd/XNQvK0aaMyVgEb1+FiFANewrbKLRxCPk+FiGQD9pjeHc4dK99HUP4kfcym2J6uffXzgJi
3RxMmO1/B2nEg+1f2o8Yo2mYV6sr1KH+DnTaS9NgFotquafiYEps65CyIx57ImVOshOc/HI13sgm
30pO2VrWKchCJ07n9jUfYv4zgMAAzBpDQzsWaxRhQ7CQj844NjdaNED0JRQx0ibiloKP99uD48SJ
E5DeCERJ6xKFEDAlyfAFJbot0uaTBJ160KJByr5Bnin1k828iU8hNZvXOXGXFJWdgJKSB5eo6smR
JvJKk+ecdBvSSvJTAIH/6oNbbgt3Ezn9IeMHAWQhVFngfqjiHcuLVYJbxmy0NxWj/gMy1y9jLUKK
RSyM9sA1zgKxPKgfa1mMwJXJkm3bP3iKYdUceYZARH7lJaqS/Buu/7HQ9twEXmv9QGlwj193cU67
M759FX/8JYF7kSmypYGG4sK3nGrfRuo0wqIp/+wQiD0wnzgtkRnJZavI6AbaAyDb+Vab52+kgvLe
2sbSMdg7aCDVTETMQIWrnR6fYlPL5YOUmdJ8kXBrLm6l7qC2CCsXYaxrKNVQoTZTRqQBVpaRxOyD
A4XpZRcURR8865Jkp3JdtOMKla94xtwzB0cqywqBaTfsWcWcVBT/cp1JOf/9jpb43/zoXL45gap5
q1ShUMAJaEt0vzotLElxF7yMBKA0g/z8a0IWgqwufUFRGGjnGOF4S3EWh6K6iM97u2zSXGs19roL
7G6qwaTOcu7/kAlrRKpVaK5tQKfNAR6ZEP2WXicfY06Mx+8TALm/FU0Q8zbW5rtWg3IZ25U5YhpC
9ko4cBdaCQnYW8vrdvPbBWG5JOQ6MvvaRb+AgZWL87tTrFG7yCqY/b5Eqb4GGz/uqZQhdYh8hvNF
FGP+9t1g7NafE8XdPpbAih0zfJfQ7gSuXB8L0ZqgCIFh8vzei2sFXY7uNCDL0+jeonIem2OOoReo
cg6b2h7sn9xb3hey6umZH1sIJ/+d9Aqbz+pv2rxwEl8hGrsjyzg89dZFEtLjBVX3mJK69v72ikr0
cPLOP5hGbUwkPsffgVZ0VegL6udVhj8ZcfsoMbnmZbTPdANjFvSsZ9+OGb6ZsHaVDNKIrcfb5ItM
G4w2NpaU+GqLVIk9jTSP92VtLCemWf89pnVnyWU04XoDgIVk+koJ+DnUKyj50bxt3jJk8L+LYY3I
f36xlfF3mIIGx8vg3Xvre3q1CisTTbAdGjKQNCAn1dj/hOXF8PotEQjSsEpBiy5SbePBuZugRtXB
FQOvpmY3w0jUioH/tr+0SfNTasp0Bv2s5AhaqzpxqkjmHwngoaQh3I5ARi9C8EWym0huu0Y5lf2D
HWzjneD0i1O+IDcsjoYso94Yoy5U3VNX4PNMHQFe7ujx9YLP/4QYk32Vj8Xou71lUhMDkKYF2dQP
wPLS9KwNROPq7nbkSPcQvJK3LMMaXpHR9/VcVzHr5HSIyN450HuRAM+56LcqjwNS/ZiCPSTpJ8UE
6kg5Wbtfq5Fv2IajaDNfNYp+AVdBIVqrOmxVWpRa/i2nkn6S1MGl4UuSRuMkgb+1usD/wGi9YMcE
FvKNtd3hgbPbbCN3m9A8Ur4pV91VXq1CKdSft7vqZ8AR+L+jo560yVfJrKwH9VdeCGtEGRI+Q2wE
VuZO273K/fmUVA2QNFS4+ytWXtCVmDCNPjKLsqhP7+dP4lmgNhQ6oWDsxco1Ff47BX7yl4Q8QwWE
aXnvzFbdtxB3itBBLbOlYvX0oRfxRiX9CvU6axnmNb1xdrlD69mSrz1y+CBG+oi7vb/NFS3EgsAd
/HC3hvfaZgFcp58cFffDmtzrZswBPXjy0jNUCzWOvg9+AEaCXJyPtyXi6O9Ibm/QMnXN5kwMAMJe
FGRijXNv8RA8xH0qqcbnavziPA2O+vNwpwxUBgPky6Xu88rCeziaMVgJIgOXu0Z2JgQ1XIrfKvWR
oh0CBC29inssW5B23zFoq6DNPns/qBcDfmdjdNDdwKrnF4nSCJNWge5eEZ95j1auYGQKkcKLvvoc
eHJcav7H6kUshyf0fKC0jZotBnnRA3g0YjDU1DaxYGYIgP/ZubuT6NsxkurpU1Pj3QFVM9SbCAAU
Xs0QYVhhNlCn7lLV3vL7Q1Kn7F+CFAjFv4T0W9bm6s4GU+X0zwRdHrcdd9CVW81dtpxyK97oKDNr
jqqrPNUt7AwiPlPMIVjWnPdE7JcjoTYWn2vzktYLpv3dJivY5TN5tRFaQxKdjalrAiTozY2k4Syq
joBBJqRMcM4mzECP/TRS2zMuIhcQJpbpJfdYE9i9K+YLyCx5p+qWLFx2/oRyYtPkGU/DvernhvvI
89uFZSzYTfndtLcKRoiOy3kR5CNZLDOOp/IAHZ23SmjwkAt2cLTMIBNu2FjuzHw7NEFyXBHvw1uX
o9pKSGKjJewnyrb2Y0ZyfnKaP1GAa6On1dKuCN0+YYRp+t8UpgfJrcTD5FEsH+Ph07oc6/JvTBuC
Rl6NwrYt9AQArE/ZJTuqaU2B4AEVsd0ZtEYdexHcuA+DLHdj+wYA4qEeJyHLGsjGuTLuWTI9HYNW
Sq6+k/debzp5WIJKtFNGbRIn40yfsjvmMlXl2VxJG9M1EVtw6GRF0vouMhXtqo9MLRCvEWnMs0aG
pwd2aeBNjeMUESuPBbTArPlkJXTzQnH4ybiCaThJ8cfGlim/eUF+xvrS3pKpGxlYAbeO9o2g97L0
NqPxnTm1RHI1HBye8HzWACiU5gaKczyvyzLC6gwlMoJJzj4DeNKoaEHGDN2ZCr696iHc79k9eYjN
5fVLVUaSn//3fGlRYFaaW/nj8jK3Bnp6veW/DgqjnYqA1uT+C4YE23ejGRY/uTOSbO9PuHW1ecw7
juhkXSTWdv+whMI7x9OYOJeAg95pFRLtN8WxQ+xpoRIBqD/hCL5rOVplV3MUOElMYe3xB/Grh7oK
u19mqRQCLu8wbk/0REALydBH9VxbxQthi772tZNagtOZyllKT5GlVNQHG06RPLfmY4CD0DxHqlk9
Fmy5F7tAWBGBO4HQuhY1v3ZHuTpWsIVMF+5bsfEs6r5jXpNuQCO/umiVfyZm+ehpRrQQBN56sXq4
HX+d6iHpAGkBg1iQgxH+NVQn4PzwtVG2J0hom27eSkGWWRLGx3Y1A98iYFId+TilP5GfMEtpMrqM
kNEbcT9wLXKiJf89Q5tzP/KmR6Yw0adbCCcqiapFFKD8GszrYjMp/uhF6iK/GcYyIOsZLc8dBcVL
8z980+j1ooLToFEGGvbb92246pdnaxC/NSzFvkLwPq5WPqMUS4N2bQ+Dg7uTrhnKfMNkh2xKwIwp
GHhkQjYwATmn1llJ8/hyiRHQPLfs4O41OIwiboFkrkAg9Fc+DbNmOe1DqWKdkBQ/xcdOiPr3/qlk
+RzRPzEH4h3oG901b3Yx8U9mAq7niT5Qxl8mYrF6TbxWjYzkCv4V5UStxwIlYziEKVFzUy5KspiK
C0zlB6UKhc3iwIkIY8Zw0Qr3cwFat40CSGcFvIAAWdesrEdJSrau8s6j9C5zEI4aeg00Kaae/ut+
thH9JsqrWBiJ6PPfhWnIOAEeQkLubCRgjy6EbQH3oKkZ3I/6BQucoYfzuTQija06iXyPG6t1x23m
K8cm2zIswDGijfX5DBpDlk/XGU+2wUtQv+nb7GYifCwkWlzM5rCak9QO8TvIO/gn8+3+l4VmJ5Pn
ec15rk8ocx65XHs8Wusg4X3PLCNew+LZxo1BeG5fo5bBruYGVVUbaMqzPvAlzbiYqXfb4U0ny26v
4UDGBuLYJ7kuTGOeutdBN6Tml/+s8ttcNk1VjKXQNWVb/ah25vORcAJ8mw+aMbR+UuUtUyVUzypH
+h9YxzwREea7NmQXiXD/LYzyCQ7dl1GN9mMpt9p8iEz1xhx8a2L49UeMjl6IYMzlWQSz0RTRj9Q+
nKSlA3ka3PFWmxwJeyGL+QXaIMyQby2iGfCjCUDr50kKG/BJVUvZMH9ALWqP/SfEtkmpro1kHWPl
BakhU9TmdThNnIpHKZ4jWqBixSd+XKBfYmmDlNChavJxnUniswEINUgtkiiWgZrYPm5Ef3JMH82G
QheNA8T3nZk3UkVpVhDlOJqIIh5wCtqUCeR1ia37/tkV6s+cqEch3nHb2+dmq6nZy8Yf/LNA6Ra3
bg5erhBAsRL4SGdUN4Qaa6Hdu0pGcrhk5mVvADMd+ropzl1m9cWWUumERR5B8ZX58o/tqNOXBCp8
IbC33Jajx0sz/jrQhRtyURNGGMlvvM1T12UKlPn2U9ZKqdmzRfvHn2CfBVss4zbmL8w5bGQ0Zejo
nHN/PEDHQ4Wk6hIdyBZ6WdLhCWwTSm7RCWpoYal6mu/dmN+hXE3HRxCkCK4TFnFDtfini9h3y+9B
eac0ziW9Th7ZdGng1JmnLLw+NI2cEVaiKlNCBT0RZkPZFC2tgG2vNHDjs1Qn5+dTO1249o2vSWCQ
FbsmknzFoGKJ6IlkRxoCH3YZ3LVOqN/sd4MYPUz8vL4iPoLmtRdf407IyoTuMG9sJgwoOzqJKVK9
XnhEsI0BhyFELYXx9P2JVxj/XdG7EKFhyqwlnbiTqTEZ/ZcAg7cQWEMipBvpBikqAPGbOm9sPK8O
kY7Qg+ugX/VXvayKp8dsPihfi7YVKhLya5wdAm/sGp/xLVmH5IcayzTDadFQZHEiFlvvLjfdYIGn
aujPbjbiVb79KzmcRguIK6lZgw+I8RGarrzKA9LQbhCwUKH2aOcjSCy9bHgkTdDQQIAtGT9Eseix
VItTBZRoOY55jDyYG8+w/X0PA/2kLj/G6st+8lmfeTK877MDt0S56+tNlip5opmHuY/hHX5ic1p1
bAtj6txVUyQf4i06MPVYmJFWrAdJRYE2ZCNLCEvkgnFR7MlyIgxDzI/Wfhn50GOoOEU+kQqZcRX0
u9jB0DEzX8R+wiBBBWYsnDh39IWtqnvd4MNYtnTmchH57yM2YPyziYjv/Tc4rHGAvk64XrNVQu8J
cMZy+MrUPocEv1/eid6yAXxDenkszQ6uNnDQa8IFZR8L9AQAfUYGSWDLoXi3+VqyUTWYIAPWtwHQ
htCQhYlGCDE5/FAmE4/UPvvsDJw9HV1F8uJbbMr8wDZ6MM7MGbY7zWR8XMNls61sjsE2JIMFgBFM
fbWWprruRrjP9bi4ypG9KoLApQ7O1EtmMrV2CwrEJuMt5JhSETQfHklE+YHoOiVg0ugaq9iMx5xC
VYcbwsupE7e0s4D3srmQghLF31uQK79g5XD30LnYWpdyuOIJO1woE7bgaEcJPhXQF9XondezPOjW
v/aYTCeQf9FyhmXXGg3h2kVa/uZ0KkNHVYfkK7uYpfo7u/5/zaY7gNh5bt6PgqtWQbsDwEj379eq
PUv5a7vKOzOGwuEhVUR32TASoaiHYv1/igGOPpivQMuViS7Lqu8ccv4F4zOLOVCiQiiwg3iPmahF
Rg0gj5rNQD16DC/YVABqVqf5i2WDDEa9cme9dJDsch2NgO02tdrBjoTrww/uM62US83U42cvV4Vq
xpTX5XMs25e2ndGLtgC8OLbaaSrGjBxtYJ3UfmfwULeBOk5nNd4uwV8G2RSfjtJG1OyOtqT4Oi+B
c3095PA7ZNAGFKrhn+e1CUAcCs54POiNa255gni2bTt5yoQRBmsQHjtlvF/3wbrwy8Sud6M6rnod
QjS9JXAVuHsFE1p0JgWFjsvCa/VUyeCLB+5WN/NLP8+/8biepBlEczrKUybI/O982SacjjcRVG15
mWrnhvdPaqvv49m/WXIphZvHUcFfhjjjSUyAi8IyDEYtPGtwjKzgXN5gJtW+mdzF5wBrdVhwn6R3
XKTkmKVafCEzCoyzcy2bV+j9INbIs/8NL8u/hfQIHSunFiZfmg3xpDGyIgcxs8VcXpZgG27nFdk1
ASTAnn0QzXIA/rYWtx5PQuM35N+M9zp8X28ha57Bd5bvDnkrME4JeX/x4H/O+XR7V1+6bZD15p5Q
QDtjjosipyuO+9RpxgFfYwnLVBvzNg0KW6jrUkZKjPb1H4TgX3hHk4DTsBWUNpz6/ppM439/VX5U
aC01So7+bazvHuW79j/duscfnLX8ZK1+0FlgJ5dhD0VXN6FTyrUYQJu8vt8pY9ldJguHpBdl7NzC
mH5RihPtbx2ntwT9L/s/kDa6ksYmpoE88x5nsMZrxDRD9+CVPsS2e87BOpG5k8G1YLj6G1mbnWGS
X0dedw5S1RVt8eog21+MhnJKdP3/xc22oQDQLLJsSlsVbh7JjZ11lMGch7EqP4JYzLv3KMz8LU6E
WbUbfIYz36pCvZq/iUHKh9hSzKEfItzpPmF47Uef6e65rrBR30hIqtyBIOIPppWaO8bmD37xpkWR
oN4zlbdw1JXm+0JW26PSyVGRflwSNBEa+K07UhBgomknb5ZMD6JIpLP33RKsTj30iqysoG8fyFmQ
tOq86kEx+ew+p9PmQ/9YUTdDzF0+1JqIW6HTdy6OI7R3ybyU//bkreQiODpT8/VQtnQDtjbkUIPS
uLpO5Q1Krz3xrljp1r6yX725Ijiqc/xCNVuMeAPB00byaibFYsbYq/YtJUr0CjJCw56HjK518Hzc
UZt//c+nGAOCqIl+dfeDt/myhJ5Wp29loSKS2wdOzuu7dFVUCGraByFAIyXkYwtUO3Qn+D3jja/P
9jBtTHUvA8R5MH/3IHXVXm4/fvif+QW2SnHk9RU3Ohjrhoe96H0bAVrGzfCwIZ7vw72Ryqm4Jwwo
fLlQhk02JWuacybTL+cxMcIJXYRxfkkjEIV4EliUO6xnKbz0tGhx2Pgojm6OYCLdnkYx2GudPYC4
JSkBU4xTYE+yrP7JaSUtEM65wmZTvBT4jC4T9X/LS7WEtgWWzg8ZJ8G8FobtioZuCTQHqJa3f2R/
mbOzFs2Ni5MJITPZHuK1e9IwocGU2Mql68LkuvNC01R9SHDh/MmocU1yDk3l6q4o9MlSxlrUvHOH
TDqI6MhVl4+psTOLYkdsDsxz4kzihS1j/M28gDGjKJIOYfpdko2WuV6HyUJtW3AzLfTVof+f61e8
viFzWbGjPPh6PTp0plBUtvcB8/Xuo8529qduPRIilGQzHO36ddp9uTQ7ulNoHay/PxhCPpKyWhLD
phNPNFbJKNte54HkUzfJTNRtB5xdmXmRb8XtfbIdOg2s9rpQ4Pst/D3Quni3gnjPOPpIAAnuVeJ9
vQZ7X2L5onfgavaiMPQlYXnK6T79BDQR7SCE/oe+B/DbdjeeMR4VLwrLP6E5CqK0usJrTuu9b/GD
d7w2/gjm6K4ijHufeddqoCkLuYSFqPexriRsYeuQlTp0jcZcA8R62gq1Jb4uQUe3PfpNorBaFQs1
2RU27DeVpZu/X7L4rXdAigPTNtD+9Gmt1aOUqm43wfC4wCRZ2GWOww/MGwx63+IAZpgcFWPiLQIF
ZJThNWCDaW+R3nPgB0U3qNdeEC0ImBz5BI8SM8niSF4HU+HGJah/VYJavFhCJFCN31C6RXO7bYR8
DlKfF48bGfTStq6uT4H9NjKrcX2FgRaf5QOf+KRZ4xVGVc9ZGe/CGYeZFyvOVM9eF7bWPnrihHHl
aQ/xgdg3YnNS189dUP14xCjRH72bNLZiz0Dd+duJNmreZj9faHiTEylmKvomide09OGR4A+7YRY4
ISNufKlb2z8olH+h/sDb7OAfyq/iAoreNEMJZWDlllvcZ7nyBcvQdHz7EqiH7oPvUWNJ+9I8mmKh
j2aGbW8muGPwzuw/0dctyZohCANeH7cJ5ELVzi7P8jtFBT+BRaUcHfNHsACOcbKG2Cg7fiXfrm78
4vnl2SRXU7beHw0+ERkb5FemKh3H4QyKryAWxFLgqKqH+jvQqCqY2BSXRQa0OAqEP+mN/rE67/Vu
2kl6m2O3Z/q29bkW0L5BaZ6HmNUC4+xvkrsSPt/r4XZfK/hKp9TYHsonNhkgeLhQ1T26M121goI9
JtFwCVM8LSvtwt7lFjJPBXjiEX+As4VI5J95oSAO7YYBfhjbcABt2ARNzApxRQZHHa8bM88JRTbi
hHJerm6SMbdsGmdYTLw/KmCicVUqeSmiVDcoI7O4lHiJZrNH5EY3Hb01sbO/eoD0tHK99Z/hF5MC
MwAhGwIHAWXpiZRiygzkrgm92CZAVAwVQu+0NHYxF1AK7vVFY1YSD7CRjhzYqvK3wP69fUJ6GfWx
oYgR9cgBLHDj0+Ij7CgDXWZrwfFKhoduLF8VBsVH4MzKNR81FZCEmBeTvvUIqSLJmjcL++mPFsRm
vJmC+f8H5Yy/taidZZ1La/2/pSOES3sT+fz3xnnnxOkfrHrJNh/nLFeRQeI0Zwpt2if7J55YUL/M
lIc3ZP2J+dyxk12AvswCuZORFpI9yd6BpsKmjiPJJukOKxLuwSKJlMILe2dFu981y9xd/TH2CRPA
SxiEh9SX82syUDBVWD3CJJIr7Awt4vDk8iOWmAWzj9X2GiWlkJZQMsMfaO2H+wpKmChs2CchL9PP
h00rPeE8v7Q2AHVTkWM0uaQSpJWGaQr4ixLkFD1CLWavI6VBlsilhSk84xAU/cYxX2w8ASAsvjkU
gCLL7t0bjSJ5nOM2cHHYlUrad6L5LUTieThODdCyWpCYsxy4XvLaEPSYf2ZM2flMXZPYiG+INBw/
a99DmSVO7yHToTmHp6Por0iBfRtQsa9V1IAZ0pViQEw/Ksn8uX0zfPX1wzRLs2bLZXqPba+hfbm3
GvQAneSIaB4uPB5hxR55Q7AtS9zmFMxKQLnZQDqhUnpefqPSJiXG/kXS8piHlQWERwGAHtUe7o14
OAtH2UkEw2tEtcIV1uo+b/Jk2GBSQDW1PZCkmnp4a+y1lssJxJ4eh6Fh36ofPzRQz4NbOwAlIgHM
IhW/Y2EPely7XvUKWcFvku5zEJVcxXAzbqz6Z7Zx+17+28QS4YkV+ovtaDKQR2mHoLjGdaOX7ExM
d+qIm8OwphGPzFLBQi0y6zWEfI1khmegYuatbYhdG29oSMtct1bzAv7az9xV0INtR7XiIzFSjQTZ
jn5Ce+r9/u2Gpx+IAHXEBCFiBiEMvChvuSzYSNt5TAmSL8LN60kthxF+VI2wz7efOhNVpsXZtY4O
XqllPmIEXX6hu1+yGu0Rf+xLqo1FgxdoDt4CDL/CsA1AExtDBzsZvyb2WGLieorO/C8VAEylmbzL
9MyDjTo1okptWadz6OfxlgU+8aLO5oF7hT0u64WsZx2HeE4Yq0fj6EyZ0JD9DoCY1VxAd+5iqPCd
FEyaWMChp8SDl/GklkXplB7g1FDn4i04PySfQv1qQyJ0WhzDwP6K2+RJelLMYRCHks+bpsc3RLkL
iIyXXXX1q0wVgO1GczF1hNRy/7M1AlCumEOV9WDO9XrFA8H8sEDobxi5D3YgygL1QWhjQogkIWf5
O5d2wY1BUQi/QluuLGYS4Wt3IHGhykbOp1R9vwr8YhGKt45x2ZsevCNiKACBz7DLel4nXPb7Gw8m
WfPlRObeRdTpWWGu8YL951Ldz2LRY7I4II4v51X6AsvOZPh63NYaBwk+47lMiw+Cv72pbv43ZQyc
6pYqUm82It7QuM7TMODyUO565iu9CNX3CKs2CinJNirXU2JWz1ZCrwNNQX1MkgkbIIq4EZuCuA+/
YUdrn9iQS5KQlk5VXO6vzBY8MK9M4pF1ZxzRJdrbHOKdopoS5MQaiE/l9uME/gNAUZ+N8qUR8+fM
j0u3aTL3HUEGHew7f706WRa9uhkfskXCAco/7e3KiBa62aux2aY0aPopi12NzC8LAuAKJXXEtY8O
U1X5zkQGpX4lFH34PEOwueb5Jp7CQVNQ+Xk2WWccTna/QwGJrEJ5bpyWVKNHhL5fECVXiKVtJGbx
fpfOpbY/sqp5Rlu2N+kdMIhscRjdRyZcK86vCeicHf+gf4phCBz/RbYVNMzwHxk3zes4xjO9BbeQ
9Bt0UM+wtgOB0F4DwYCEFgA/F5+kTozdNguXDPfQ3cYg0pnrSbQSPjKvUFApnbbLwl6AOXy3UNPI
2m0n/iOsj7EP9noE0CuKq+x6E6+h0s6IZD/6yLZQkpZiWwghyzkfev8v/12KdN9vBc/90U2jhIfN
KD2n1mc3IiLAqLiXG9FD4WbfNW/WdRgo8kvcFtGK05i+2C735ELFpjL+e7+peK4mtwdNF93Ba/px
lJyaFiSqjF3ngZ1g9oStSQd4taFgDi8/LBjwTH40/u/n+KOUh8U5Mt3ETRd/wqkJk8almTcbCV75
x70xHo0UbZvKZYwecQ3z/Bk/iABTym+GyUieGRhrb1OKLJFSF+6nm2fenjanZ5OL6L+bQ5O4YkvH
/iFGwpoFAQ1VBGk3BcgTPMfOOfcZrUp4IGs0qaoXg90V+DuJ42uQcNaCP5SXfRlyjLWqa1UK/jTk
Mp4KAL4zZ1QJUFQ7rTlgqMtK7+keLnkKgS3sqLqCfMzZjPoJMFKtXdiQoRE5VVT5R9svmxdYg+RJ
Fmm7Le6ORO4ZxPUBDK6KgXg0uW6B7Pe6OR/6yu8y2SKm2us/ZmLLWQQLLcO/UV7TQu2xf5bu3W1F
m4u4IfMpSA87LXQqCqCcOGIGf6svjlWdcv2LR9IrwBixffptzD5cNR2H56QvIyDw6NZKwI4ui6RV
wpiJIEyAhuZL1hh6N6mSkrilL3lgaF/vU9r0PNEqJOmx1f0TY9WHW3BQT8EjhMpwVEGz12i0w/2k
RMuaje5E8ioYQV264mMe0UeL/nIZ6OAsTh59xkAD9R7yGCkXWTbLlrw8OmEX/qKsNLF0MerYhnC/
V0SeRMqnRelCpi1OBe8DKzoGl5qiD1f6EYuV4a29PvISHicHw5VPZnWpY5Yj6MXo3pdVHxb5y2kD
xDpDSS0MUsjKBOzj4QwRhpSAEyb2IYYHRCC4cBgOEXQVG71hhCUlhCiUpd1h18jrt9jFoj7WDz3z
quK+jOoNLbD+Kud1g00x9kD8Gn+vO6il2ZcqiXHwegOM6nJPgHqgG8d9xyONO6wB9A8/HSxRN2Zs
fPNYtVOcb6H9mLRRKYUiNr7izhtK4ExrKg+aWFPC171tNvRrvH6Cem1MqHNzux3N904FSW8wbYr7
HDih2NrLre6/B6LF6OmHS7uDzD4yYeihYD1gPKwQpGQMUBWweAL+ZItjfUwb0FLECljKE7nz2IZn
hqvL5Oaot4XvIh3cfKH35PLQcMG823eIRlf5HLNFmMcIJajfsEjmm0ldy90NIMiD4S/UMdb9pXsb
DYc6YJifaEC8P7ykASC4wsSAWxJfta3zYare8+ukQHtd9m0thfgbFR092raJybyg8eIwBJUDrHY6
eokIRF2TTnHXwU7SzrTot+0Bz8JM5RvJrBfcOPacg/lnGy3mB85nrmeWivgdHGcpsQ69bjIUUDCc
2NkSy+sxFk+1gzZ5hn+Gv4xSFxhshOQrOOqc34bNEEq0L4vHsoTZXMVfXd/PaXNK8Du0VJNR6xvN
MxaOwm7LhC1gJe4pwp/WcfU86gLuDqb8+q8vJqX1FUbsnr/eOEJiYptjrxTI/O61SDLNgGrXydTE
Ji79LMHo8k/4zXcATsZrUCyzv7xCt3T6NzeOSZWr0zIq3bQ9CJoYNuMIujC3gS9EUB+GYtEnGlDf
XsiXR/37g2jI4jQ6cTDkZSbkRqt9jYVU+YN3EBdret9kDGgfUksa5mgCSQs0cyb/aw/CKjAEsgJG
+CrfErxAB6eLZQdSl7ObAl5ymMet5SzcIVvb0Q4B6vHkThbJuN87xxA7D/ZlRpK7uHGWfMbxae9P
CNCZabp3RbqWNGzVscYS6NMdo8scjU+EKvyL0ne3NIWwClqMoFpHpsCR1dVl7n1DcMaG4rVRp9tp
BHJiBLordrAEQ+MpCDUeHZaOfemnJsHkiXrqOSdixWN65oferj3uc4xnKl+ekK7MZuUruYDVRBGy
EySJFClGWp1y3bsneOtXeRgji3BIoJRJleiSb4W9QP/+6D5pcPW63E9UPdo61+XpS8M8mlEltbNW
GSdhfTCWbtubAybX3LYpvYC7uTS6EP6nYxwwVAnROTN6G8EHNO/QskQG5MwggXdgxN8dmBngl7Ri
WeKeQWggqgX/Wv3+00RV5bahdZ5xu9RiQmWdrR5CpZgaUoqvkt3MSWfjg8kvRU/ufbBnDSduXPdq
ETaa7AXtsYIziVkc7n9dNqJPOjHuzDrcCkqtKPLNGNjOQObL4a16pQpjOFrUIyV6xNR7jbVIJyNl
uIKDM8zOYV3JtGNAjM72LxcxlixY7pUadFVSzn/qg+jfinTcvbNmZSN3qSG6KThbgyiTrFPPyofe
xWkVEQ/3oQ9TgfnciASRh1q1Y3zKlxS3gueGMI9vY1Q9CetQikdqLZZTL+otLSldxWTeAMFp2zIR
iuXhdCUBNqRiQ+Tj6X0+Jf2bBp7gdixM0qkrTSGiD+6ZBJVlAmi7lZfpb3sFpcLGxgqHcFypuP/a
jzJwfkNu7gBTTNta8l6AruAugB5ZMCl4LVrkWTKokTpEioKhSeQm7NGMqZau+aiqSxUgz3Q5QTZz
JXnxma3hTPdKbL3MKQ4UbrMG5xGaYWsy9vzyOh9f2asyLLkFdwcHQulwgSfsZrMBrYRvBcS51o1F
S6LuorlqmChvwm3zpvs/mQiFwgxqOkTxnpRAwDoycW0rNZP05rhVplZM9o2jusS68PWDCEnsGRdr
NXHvPdyPtYCkeOCKd84APyUnxrNgmr5hXlzp5n6X7NpsK1OJ9PV7p2Qt2SxUyxYSKUhN8V8rfPlq
G8p6WAvzphPwJ75X1z1BZZoJ/T6vhshs1Pewj+HQFYoSHr86vvMMv84bmpbAoefZek8PWcUOSaic
doKg4yTKlNUpsqbfLeRN+8gawkheIVq3QxkTFr8VuxtAeb0BZJGMJzL5pz43whDxhseZQ3neUshF
lQUqC2N+IsGHrbhiKdluL8DmMJOwBBga+dhT6gaHUGy/YeDIzSSQ6m7E309icLoj9dxFJ2z0eYJS
R8iNJpblvdjINn8No9rMdmz3XLeFxixautrczPmA9fI16yky33bXt7XgmFD5CJV9ZN5b8gh98V+7
tcXWwXf2sNdoddaqeFfN8YakmFIuq9aA1ZHAxLAPWXnUBg4aFAI20EmceIO55KSHHgMCxHEzj9Ru
XTgdFLz3pu/s09t3DHW8GxxCDnhhJsNLUcJvG41zDkE/e+Or0XgH3S55Ech5iTU54eNV8/anUeVj
G1Qzij0coia7me1TGOFitNh1SVwmTwyto22fgX51pVG6zM+Lpz2fkR+/ypAL1Sd5+SNSZ6XPYSjc
8pytOHWjU0TPcsSTspLnrbWB3s6wvPeQ5hAKPCIpN3zBULxtOUhcEPVhBWi4EaSPrNj0pknhNhwl
9Tqppmtx2djtimvxUoKRXO6ow2hLvrrmXCpcqdN/MPIc/PdRWJq6dunekN+ekZQkG2qO1i+d6SV9
VMV6rWPkZr8TvaiYnTKoCJCMr95cSrR/2mVBR8lqqC/fQI33HEsZGBcBSGT9ic4K4LPHUY+wawO6
gy5FWdmchy8mqz/PPsMor8AKkLuMUwFZJNnCw3//9bki3Sv2P9peeLBcpkgNwSlDwi5Xkp2s6J+V
+6aHJE/TZaP6Pz+b8FiUW0jAXAr9ZTR1Y3XLI2LJz3bzDf0zybEmusSDC/6qswwZ6Sxy8rsznCqT
GlJT/pPe1BUVy97qUmHm2gTaZ1SuTJ5Cm7WZmswrRDLHyxsBP4CwJh5xQsyVoNc/UGNJVhRgF1ZH
zQ4GtrTqhhpiYvBxjM3k1GgcxUgp93snlYlUi6ajJ/UBmD32pv+G+dbjIh1hU/Qzlbbfn1bWfnfj
/aDW6Eg81/F1lnaCLyfSq8BADm/gD5eAzMgDstfRXmotBq1KGIviQm0xosKVnNf4KFPderbsnxou
gyEios6YHpYn7cQ9P3lnxBxlzg+31DFp0cHzwOiuwhzYpWpRMOHCtM2wh4zGCpFkJtkUHZP/6XZX
m52tPNdaDJakvP5avnotBBdcXJooCsFAC+zweQ3ZQBJCCtFxM5daCqksPfjA5EoOQbAdrl9CWUp0
6Rju3xlugTCdrzVKuDZO1B9Hjoe/gC8vjCOf9EzB/5Kk9P3AR41jU5rHZpPP8qRCmyqmR7woJyhB
j+8C69h572ZpKlSH++R6fUB8Wkt9YbanXXZj/BjO7eJA0OuDTCmh1E2AZ7saSvv1O1hT9ZtWXLEe
M1OioUIffriS3sdrb2gsQDNbmW0gs/BmjD3cU63zzvGbzprHV5Y5KhtTQu8XSkApc79rc7YemBrd
3tVMe1xQBSuqvPLH1jPZMflA0aEQVGgfc5NMO8trcQiYLTHphJ93B8yUsSNVXheFieZIULClXoP4
8l4QdwBmnjK2Vz1l4ZIS6w0DtxMymRJ2dRdnQ2I4VERfhh5Tzf96NsdxecHsy8uW4A7DqUHWf56q
qDe+WirWoqIgCuj6JcHsIGCc+gjcrdavOXclqJF22l7224OmtL1p9eA4+5GzOmXRpIRvd9UE7uzN
0ghlOLnnij3ZyEf28a6j7jzb9io6IcVj8hnoNFf11gFkzOVTe7s0jM9u08frGrVUuc4asb7/T8jt
UHJQ33gZRL7R07+DmaU7BvYpNi3YcKn49smDo57GoXEXvA7AjSeF/4ZL579cpFh7aAMS1BeUSdK9
0H0ysPfjlkV0rjXXfDzf4H9SDb3HPB9c0DPnwWT0IiCKuNntGalUo7TrMxI+BPEcEp8+DiJRrmbG
cYZIApqZT7ixd7kcNolqaQadAeR0qqEkBAGvSrEi0vEIVJxt/tNIjL+iLHommyIZJOjy6swf6H6X
yjoTugbypir/QR7zMG/xZTxAYHRT7dVed/H863/DVUhk9OLN409A9BCApt6uUFmfo6qxSILbS2VX
DWbPQlGFRikscYQy8/sla6zKK0AUD1V7NwzMgfInEIh3YvoGps4HzM8D5FG/LJElohjkCUHLMTz8
IavnOKY6yZUodKtxlRWYKlsnun4G08z18dfsdehBB/HTWgQAWLTc6QM6zweM+PfrC+KBm/o7uxLl
h0bDwAgLYhrqAkaqtwlxZIYMXDZa28/vbu/uK7YNlnEBVsS13bj5enVfayLft9LBbsaguN38HPza
bQOoMpc9lnlWvogPZQwG8jCagRDZRvE2Wyvpq5N1q6S+m3ukhLXB5Nj3mmhVE6YLsiEgkiFSjnN6
J/0JpZwZamRsIERDdm7NAqI2+PJV45+3mUVSypbpQIJRCtoIf0kJV+sllZQHCZKIyTfTEtrrSebw
OPh27vhfobfuLnmMR1DEZ3CQxDjoaqBMVGFwLhRj5oGKczIY84gXED13wDy7lAiJUronTcsB642B
T4lG9tX/GetbpVPfEqUf+HBfnol7XiOvJdW5Qhnir+gzha4iGDqbWNUlhaj0uJUzmffubAANav1F
9k9yaZctxoqZd8lToBDh8wGGG4taXz4hZ1Zvl8ac55C1DnsV2uOLPU3QeTQXX4zGn5vBB15AvBza
laEgfNO+ZNk16u+AFO9sspQMBKegdmCZEFV9zPconVB9wKK5e1McvOdB4cybZi4wnMP5uNp+Bfke
iUeBlcMLLO19FtT/mBBsBchDKfX2X+bsGZaxClibRTMFQIfLSq5vhINlG1/3+4ZFzj5J3E/R68Jj
s6RmxCRdZWqHdJsXwrp1+vDiTNl5D64vMXSO4Vc8HzmmBvGLMeoz7i7DK19Z2DWmmVIuCH7/Lo8t
qMPC3zTywbyinE/XOFNFxy1HJ+c18eSruhn69bd8Qf23PWzVsGcw/M2B6r8rCEMc8RAVMGE+ZUp2
JB021I+2LUfY4jMNSv7v6x6rWDYJxNP1Si/wANkSjdKOuV7UOdEUH2n6gRjKEsIbUPPMzJ+c/k4R
yBjhVfyra1/uE8g9yhrPjDER28e/Cv+838Nt2EltdWK9x0R7sUx4zYNoIaHEraAsDcr4lnNCxotM
4xUHXC0bnFAS2qIHr8MRMLY6Eu8upA5DCtWCPHVEXXh4QNbYxQqqBkGMF/jn6JodkiTRLaaCPMAH
ySUmO8MThURoFrYbOvC2jly0Xvxx4kH4VV1SnoCkQbjlGLpgoymUPlScMSTXmiBlL/nNEQRnFsOk
jokHtGxT9kK9nvP5BUlszz2gD/FQkh6jWxlMnN94KemLwJyP4mfePBM9mFMllyCZgd9Lg7CaAbHI
KJeI4dsjJmkRHajOb0WguaFkBhz57lJz7dOTHzxpoQMKNrS54YstvkFAvSV5GqpLq8WHfj7K2CN9
/PcpwRbd0nKo+L2M7QPVP0O6D5f2sJMANujITeygQCSM8lQM5exG4OM+B2uwA2f8yqwf0a2WOYd5
PxfrZLutIHUAdAE9sVTGig8G6K7BoD4ocjpxCD4HL7p+3I1JHYLjs+5aS3aexnRIHO/YPML/4xVR
dceMXI2cYvxYasygdm9Ovsl73qG2f5oOJvJPXsEOEazJxdnZHvtGPQvsqwm993TKs4hsXHmLaA7H
yP1Eq28pAvuxrBUsL8E4PKkOFdb/ESq9nodIkq/L1uabOe62Qnavkh48o+HvraS0QpzqmT0x265U
9sHY8RktYAn8PIsnCTMyxd3prjSGRYa1O84IS8bcMd2zkTHngvkGwSXLD1cvirhz6U5liwF0qXbu
DL7kOcwknqf27SKtsxrdawSRDUCaasbYoNpRyjuUqYNvnffNQgKBragVLI4xDwuVxTKPbUykgue3
aj2QClZdVf3wai5f+OfZEDFptKYg/B3r55j/XM2zcRQyrZpQnJ1lSNLDCYv5KB1NX3zkoni6TWdO
yYjZCI6MQQITus4K8lgwhZ7FAONcH2sPyn6kWXrkP0JtK/iVK/E83O8pYGE5QJ7O8FPw53o6Hwr7
7n+v8ms5BphhtkjpEKinRDR36HIUOGAMVf+9SgtVscZ7bEjvBcs/BWprP75Y8oZJDeIUqK6Y/eGy
TLiYVtUhnvMBwqM481W1O+SA7ZXvMyuV6jnhoLok3iuUhz6bJZE1F8/AjBKrJ9pQ5qpdbfGHqTf3
l7m4Q1f6gxJ8EYLKeJ2CK/GEDSPedfJo6PAvQoapdqlfiWU6Rkd3GVJwAeDOOUl4CA5UhFRuYiYS
ZRJEPQMMVek2O1e6r1EgPCV28HxI1TK/E7/Hvkk1wk4fzi3j3MlmmQcmcLqSO4USHYb7HYpICbeW
tnEmv/J9VmXK5XpKjI7sBMMIrWkVDXwKdcOkt4yxx+LWz8F/ssdHyYot4bLhzzFcVtmIvsNQbi25
0AsgDdAQZGApZlX8YBRj2cFFplgWKNyHb2o4LYIFO1zc9PFtM3qxJ8g7POVzqjnmwmBhVFi7zyow
nhR24KLdJ2UBuVX3ks/liL3esfQ9Kz7P7+awMnWCjti8aaOoirv2951tzPwgXW/r+AXXQRs1MhUO
XUca661sQC4b9zDbuDy9gZ1ZnMgyTUTDbHoeHbIsrQrt9PQyyNZwZzFHGKEUKvvN2ZUrydiIqYqz
0cSKMWNNmh4UnhFd81T7jXBqc6UkPRYVhOAebv5f2ntc7asJVh8v7PUbh659bftcFO4vscQsTXfU
iy/EEJivTEGNXFcnTMQwfA+LZ9+uZ7FvzqRm94/UGfnIdEwo4UpVKZZrP0AECpk4Z9JYxjAVFr6r
uEhr/7EP88XeSIucfvFeyyYaJITRayNxCgojyGJE7yvrAikyMP7SuC+L30jkCXFThpseVHkDdRCD
aHrTm7zbjlCyvwwRM+m/gjl/X7PH9LMiFB31Vkbe9iyPYUQtfFAmsZKWR+DsFPxVK84nQITY+te5
dUPA7C8sGTNMVRn+FDRXlTXxO3geS5WqqCDH17DNgxZ0ZPQ3pQVn2Ff2gpR2T0odlPLcCtehfqDv
oOUxClTAGwx0RvT9uDKY11G2ARO0tO5ptmW0/DZ4HeQFYU9dsED0cpgtWVTFkfndV8hNfSCvD3m7
MFWa2O5+2ps0mgeFgcgrpPHfFXzZA8qvt8R2b5kmnNM6HZGozTZsM1jkKoY+b/HbTzG3hPr6RVzJ
Czi1g6LB7sJ1rCmzHU4dGwMOExAQ93jiE9NDhWOGsHOxNosPy6eHPuJg8rd8YRqurh2rQftBRshf
3cFYFxyoFP3YEzjdiLNdZ5CFMBqSBQMC1/SnSGA1Zy/EZYKKAGFBU4tu4lQzzl+IuF70197TTkQY
xupF15sClDj6uWyF56OYtvCmgqKftjXgy+rjbvMcMOav957s2Y0ljxrJd5lScr8BGMoIesqJzbJW
ifV/WYhYNrcjRax+0cCGtehsqdfRs09YL56GDn9k076zQbDFMaBz58iwJJd1Yqs/X5mTUpoH7bF6
aytU7RcltpIzs343MLBMffBaYWrOKYMwgdgCgfbuPyVHDhK91biLe38xg5fBKjDWz3yRyXeJRxFo
A6nY/1O+4AcIzGBEDlmIZ2PTSQRp0jGR9hRmx2sLsOVZES6RQ0OiBOtnhaAPu1nNMYjYzyBtJMaF
C/vDy/GWD/9tDgP7gWrLnCEeLx8V/he2P5rgpARl0wsLCl4K42FDll5Il7oguIlXXJd3LomBoy1d
QLtNV8EVYJJOube7Wub39Tvc1qXTbOxgRMKCEFvI4qQ6c47+XKLZ3rKpPkDwLaEod20vYaDtTMnb
lYZl2ag2yw5xmNENGEVr96QKqX/9GRN9Hbm+OhhQju12wg86xbpBvYez1LBt0eAEf5sn8p5ODBaR
8bFN1pzkpIDUkzI0cL+x+TAiMD3fyqv2K1fsm16IvoSJWmLd5T6b46Vw+1xKXvTd1z9Ljkw2d8+I
KEZoXJDPFkALd/R79mscK93ZJkUnkzJ+Dy2NQhiDVKZL6fgn8Hn2fPbzqwyjatn+Zbq8bDYHeLH6
8hQc3rn13KJpJtlZnxcS7aiTBH1PXA0Ml2v5m7a4vfm7GKhdjOGR7RmwrvE9XZL7zWK6Xjaj8Hco
i4b2SKBZfHqujWpF0qm2zW1eV5tJVzDmBueTAH+NWNuFA9kus0zidHarnvC4JpNmiELrgWvQ9dED
8RF9EYO3h22YSua6fT+BoQo+VjOFPRCZIEHh0Chnn2n2LRqdRxFTZKVaAFVkyxnc/sAIduUFj/YH
ywhQfXGXWAbPBOfAShFwHdHMfOFsekCw8QjF+C3nhCYNoBm16VtHdgT272qSzi/znNx62lJblike
1UR1MLDrg9ffRSyOJW58rcom1LykvDvLjF2OFvGRgHAMa9jPW0VQP4CT+xSfhIOJN+bUKSVaPxze
3TCDIx9TCW1SakKioy17o3sO5Wh5C6vCpwV9eNP/pcpOBf/M1T8qWqhn2nw/5FdZO3nj/t7uoPx/
gmyn3QXQ8O7oQceeGJtR6RC8YwmzVGZBxD3Ih8OWYpdmJxwatPIKLKgpXYTdcJKGOst2qOYOcAf3
fhPKsDE5cVtmFP1s0MywvJ3zEycjmoJPQ6vjdKpvYRuSh7FQaenr6pu3x+fsKQA4UW0MyTlek/TX
d17DlYTw+POrP9Z7238al77ItKQlBYX6RCfePxm8z41YkU8U0WS87AltUpVjobQ18Zff3PutzzOi
QdDC4Le+s3X8dcZ/iLksosrlZWQiFzhmOFnju1oBd1ZIs6r+HvctY1EYcRwdFV1pT00B5CiGMdoi
LQZWUgu9xMd/cFnBPUCq0P84CJjkTvMX10SnSVjeXDOf3p2TjQTx8X7h6psGJBbroBjMc7A9drGm
Ns7Y49cXVqn3gB75VTnDNEfxLmTPjbSV5LCLlOfreX00Qxo7h2O/2vxKg+gU6r3V7xwAFJvXl+Rf
NS2rTylZMxcZ6rJySRoWYssa+ExbVQmUgasFbUEsfKm2xh6jhbHm/v/eAAmOVxIVkomxM9plbpkW
tek5kvcgw8zUVa0DXmat/gfgzqbC9bQfRVh7uaYOI7rEnX2jAvREs1fTRLe8XND3/wvgFDEQosJy
rk6mpjDGNkwhb9FMqkCxZxLxWElLssMa83+hw9kZU3LGCWeb4n0GvWnQFw+qFVowDqymVXP7PArq
Ljhy+RrhTtWy9x89SsO5pI2vNDWikTF9DdjxJoGvuUBjWopVuELP4QmG19rHmnKs9pLZcc5iTuBU
0gefapRBwGpxU0t5wojBSsoMcJKAbFMfKeJhRRGTFRM5FggrN3cnT+QJIIF70HobaSJA+6i44VK+
o7f3Or/WDvgslwaa4/YZ6hKYGIr7mJXIOU9m9FqD4DBPZhT1L48aAtcVZDGVEHWbP/siUUVEbxds
Lk3RY0ov1gKnyrvO4bB0Clbe32wjoC9UAaAVa3THpnZDKb838rv01gQpGqbwIQGCn/t3tjDc4csp
iq/G4mbplUEUfvFCtm+i3lsbQcbQAsQIf8RMMSpT7f+RK1SWY/w5HxFX8o+EqDQ1dOAg4424bFCM
dgabsIHWK+hmrNfcbsgmK3o+zDSZlFG2P7drPbPwaUk1f9n/S476LLGemMyW5aDGY7wW7qsene2t
dVI+7kQlr6NAgpNeQ+ANd53VXnvN5Gmyd7IdaHMmChQ7K+ygC+o215lV6M+TS6pWTT4ysKf7rYO9
CD+FcBMzrKEmYMqXWtzrCtmnfuewMRw4L8ZjXGHwc3LaKz815kSlnAeGNcFaqdhqFHluIRpYIF/I
PSMwNEci9t81jTv79xmkigDTmQ9MEA8UpUWZNWnDu7+3Yidk6tQhbOSt90I2Y6ah4cmHerbyphly
4hiIAfJ4dm0ZvS6bx+CQkmo5AgOFMb+vqYKLA1r9gYLtJDHVtDrlD95Uzus3SthXM8w2pyNmW9aj
jz82/0Y2nadjfzDbrjVTdv1r+5zzkBeg18piuYPAzfpw8HbITG/5mVJo4Ee4y8bwAXLrFObuK0/v
uDvy1bEjSaa8lRiMfjfKkWhLjkvxpLvSshsC02Wue5iBqfbdV3WMembIGulmzNOvimSH1pKTfTrv
p5rouC10dToOeAt/YCXzRw0B8IWJ4ymlm1iyx01Z1wF5U9pBt1FZTExt4eBRSdbdin7zfZ3uZpcW
xAWIOkYFNtQm2nDStQ0lZrXMaCc0C8z3YwSueNv11kRxBeB3xms7M0OUVFu7dR9UipPcR61hW6oR
aefW8sp8gtwRMq/PVzvOwlCkXXSnHlVGRxxN97EjlJnwGQYYnf5wPH116GoSBUXeh9Zd/I76jesJ
nrkc0/nZlu1M0uZqjAenWmx4D5jAeC8zHiTVHB15OghOnZlVzoV+rIpGEJOLdbLH2MhfvECId21+
7uAapao4sJ3F8NfMuduUVZ2SmMgJGX2LN0iQKn8iH4dm91drrqpbtd2lnD+6ED7FWMbEs5/gegTX
SQqFg5tOqQUWnKMOFvw77nrD6qnOmswyfEkbwLcesqAVAd5rV7Ax8QRnlPX1zLDwLasi+Cka/Vta
hUJitYn4FkY1NI44tQ0PQjzIC28WNLRRuaSmWK18E/0mZPNbql0hhevC0UPuBFkHJlRIsPcFvyr7
7kqpSOheRKzsWQnocAYss3n3wJm06oh7kD0QFaNIOmCr+ce6d6xqr/B5R+Z8o5Grt3PzllgkPZKK
sBJSE1QuwP0qIMpho5BdY0gtffA4i9AHmEvq136sNb0UflLm01pal2vzt/DM6jNKjMRKf9SOD9yA
XhntM5CmjVluzk3DxNONhuXleYkpUGok0zHJqxjalp80POZXyImfyWLkbBxwunDu+z9TBDrbbmin
p2aIWiGNuUiiwFjq971MUEZYoCiyBOyi6Q/407WnxlswiN1OXRru3MatQOsD/r/0icWPz/++Khgy
HaS9CjOtlFy5S7PZhxBAvXrcY/2O65BYPt3xeZBWHycOcArY3rglbWS39V2YOq0xSSR12shD7uRo
1RvhAoTrdgeeifHVOoePwDQs9CKdIl2cndRi6k/Hz7BULStemo1hQMkjV57zpmE9skJEFdoKwXxe
IcNdAw2AZV6l2pWz6SEWyxo/Wi2kgX9nBupW82om3n2zwWs7B1VOkOn/qapGZkVGqty1SJKfLD8j
NR8LhUUrx+0XTLEcY3z+GzlcVGvWA/DDqmzCwkfp8ZmNdccaoQxwFeNePrxvBlCstvKJ461vULtj
7icRguIMMqZpuRbOpQfOkcjbm2yWL+pJd0hlN+FGY1AC7cJ+gsAnxKSYv5DfKExuMMIw6ZgW+p9p
xJH5F17GNR8Eytwg4dqQLJaNxPpkTs98yaSrTcekTwBun4tWsHCQ7wVvFAwPgszfFyOUyBBUfhrY
7jhaucXaLqpbfKm3fUnR9/ihXbexxj+UIv7FEL8Id0K4UojnDqfizcMX6F/i7qYenY5gJOr+DI4U
7ZKRhRjnt8yuB3B5r1TtwjIFYUsnLLLAwjPUqv0hlKgVosHiUS9JLb6v5vT4XSJ3GsT9HWUMtfdb
a6TOsEnsJgBcUjy2xv6FKmduSUTSaJZfmUqspvotriLnem8uzDlO8YUQxEoUUd1CIbW5uAeImmUM
20OEKBEvKJ5EKW1pRdcLcWfCTMGP4iOvI7+JmD6ARvq9IYof/Wg5l/4caManqM6XebVmcV6BBAal
IReAnK8HNAehW+oXFUKsqM0YLEqUkybki4Z4zSAatlvZu4gSjmHJByzghBBre1Z0VGwaIU+reYf9
9s5JINjp/zSSMLcr65TkS0bWdsv1ofNSx7W/9Y0EaHBWCsEb+5mmrGerTz5zSrLn9M29nxMOLDSU
CGKIfIfuIIRkmY+Tw5BLT2Ty4FnpHRFqDBd9wwD0vyw8+7iKZmSqkoBcBW/OTu9MyexZdlAV0pHt
5fzmKFnynHIBp2fWAgRjvX4bJegORc3nblMzrR2EgEbyboeSE7Od6Q4iDMV7bTmiyyCuycfq27Be
4jOg0L7li9zbM57XYVH/VHmDI5Ymh3WrmtxutQoev/UTgc11P8BYrzER+g2UJ9f0/eIydHyMR+cV
GEiuwxktULL3HTpmS5ysptdVX/K3E5+xVPNNSQhtoixD2v/BYNoHZ8OwLkPM2xvwcLCXIczbNsRU
5pziIgWVTQwAkRQPPbdbby8QxNfAHcOuxYA+nEgOySmM2R5YzZW+E67r+FdDL0wi67Y+b+JcGM6/
hKGwu1WRsvPxnsYkrDdZXdGCPkNZPmh/0fjaU+asJ7AOu1bGpafb0SoY9NeIavUStjX/zjUcu0Ub
awm0RS+ryKK6yxEXbShG9DaXwY5HQ02o+ZlOmuv0NsrHzA9oUWDocA4wV1huWta4yWDQ7zyMwffz
SuwEU19Q1Rzht69C6eujFH45pcsyAQXJFQKv54DjExYvo1C8Wu/hUcQdY5wv/kfPyB/ub92XzpJ/
qDx63ixEngHBBS5nPZZblm5n/7vFTy31vE7BRTCmiEbI2V99hGoPPbPY5pQR+DCmThn2BNwiPyyU
iEFqHWC+1Bj5AuTvB3/diA/Wujcq1zqKUJNlbFDpG2bCm+Ux/ZlayRgmbhtxGSRH94Y9nhKP9Skl
4nG4wBpLXYFBYFAjmd+HQJgvf2e3VvIJy2Z2+5f7BvfOXFizXPMHaIGoXBSiCyhkWNC48bm0quZO
Q3+UvQVoGHirnRycsl/KJFVod6Zc3A8UbQDaLUUaUrin4uKV0vkIkkWvU++WVu4E6RbOf09v5jjH
vjJzqFs7ZGA4F9X9lQvWrtyO/59yW/eKJpjDkia+I0NWD7itslg3+rzU+mNWwx4wOtusJv/92SMb
hjs+NoEPKcR18awL7Ei+sIPrPaouw9heewzwdfWT/DCKQEQTIa6qsCjGhXLdn0jTc1dIIzrYY1ZK
lxWbH+NpBLHLPqmdsSMTf+DIgabZLfgKtHMvarK9+9oD7F2bpgigDuR4Ds+ZhRlAUe/qTtn9sKeu
66DWqCRMU3TK9uBGLQqG0iJamkeO7apX5spe7ZCx3mv1S5vSnXZ5TK61F1JYDtzXFaC7gsrf7IeU
mSHeZKDwkp9PhsYZHcptTNPhs9h7s/6f2tBJCLU3jbzr14C/g20dfKOyQLg/JMZOtOeN/yZlWyf4
8je1v60wAiSutfghzjncNtU6VPOWPs7GrDHEj9pVmDOujPDaRb4P0WTZo1u1/MChT0P+CWXAm5fZ
2grt6Xlv5usB5jjcRMBmjPJmskhq+p5SI6zQkyHX8J2lTL1hT3S+v8Wnw51vnJbfyfK3Xf6jmKUV
73JMgN55nvYOanzexMYgYwlnogWgdV4LSbHsyn+5mKfdzDukCCSnmN7IX6LMnWUtkwFPSiXuQmGF
c976HRrju8IIbDSSXPvDMuN1G+2ssorULfJgmSz40I/SpzjxJ05Y8DK9Uruuau48RgdAuiqRjPyF
4euwF/GoxgkMOBfbMzh3EOGSnbFbX1zh8qQ8hINDcClKjjuV4o5b+48LUD5rQOR/k48EYz0H4fy4
py+njfDZ/WxW7v9/ZmyEk11SJa72t1tgOynecz9MJYuEUlf0SbKqSnftDUfWJ54EsKabgwYmbSrX
MeF2YQDVUVFpj9i73pDHWdn3lN6R63GNH34SGbcjerPk6eFb2H+ZifsPPGkaI48AyhA4Cm43aspm
Q+GofDObaADdRQZgSyHijzNIRiiWml3c/8v3k8DS2H/sc1k2CFwDY/XTAwwUrRfFEKnYGVZ03n+m
FYfxtb/Q6kGjlUPiYiNiKSBZSmYRBpDNrEdm7rN3DAx+Wesju7ZYzP0M9c6ecxoKLRnbkMc/oHYY
nUf7SwmbBsctYt+heQRDXQKFm45zGGuovbzVtT4wSdqkmgRq9sfZPXO9zh5bfWu0gRj0VLPtnPiq
8jygaHqAPt1gErX7PyxzGO8YbP4n32lab9y46EMtQuz/n5OXHko8YJiKf9XdSNU9TvsYF7jjKYf1
ucygASJoPRffvznV5Ux2z4/AO3F53L0GmqFirHDR6uSoZEcAWCrOFl304sFwIjRmcEwAuY/dYYXY
1iXr5gtoVczZ7YcT4UP7a8iCERZ6VpydEV7AQKNWpS8z4Y6Yq4zWqkBtc95Jk98uR7SjfD34w8qa
NZ/CJN5UhwFfVPChYSomcX4i6hAZbfSJkc5vTgyLdSkpnWiK5E+iWXw1XVZxjHAyjhf3sFca5xgv
AUc2YHH/gpuZfmljarrDpfZhHCYq3zrsuVin1DvzP9WDmS/Hd3yPgl47r+rC8LQkG0QMiG8XPX1o
Rx/aBlvObobtf27l14eDPy9kW07kjOm13VLLdpZRdosMlV85Nv9dcs5t5urkwgZuSQKQ9ZJVOFkT
nAMAgh381RGChBNDRgoazblDndOfB7k+Xshpkn/6fK9EKr1twunLOMBhbm0uJcx9wuxE/b60Ywjh
74bUcjJX4+SXi/yhu6qM5aT4El5CCql9LQPAWow7PBDUYfKKpKwsRmJUY/n8eC+VLOCp+osgo1wD
6EEq3lkWqzePdczZuulnrs0E1ERjeqAYETiPuVZIID/Ilq7Am+OtjlImGCIEPudO86MWzH49jFFe
mvSDlW0o4w/eS3AnJUaeFwuSEhGaYuQNglTBsY7CjK32f9ff1GXyb7PFewbMlKTC522QyNlv7kgY
xgydqfBMtryWfO1SdyQg33AQU4oJro8ndZ70IOiUNFxE4dnkBGg+3y5Gp8ip5Na3g2I8Mqt3YGN3
MlSaHlMLN+PzNFOD1aqbUqusbOdEcUoT+p5fJAxP7UiXJoMXXEMpRa2bYhnmxT55o1+Z4Ejx99RQ
u6MyoTbPN2uc7BTdEgUq3sSJEZD7UFeUq16uGCRi/mFZjQasMXJ9SVWEJkWThd/wBEpW1crIu8CO
NLWA1EPkMztDeiJOkIqGGS1fTmeh9rgDUICTpjHoZsV8QPg6NYEe/UHPdqVtmKbcPAM6EP4mbGMl
YvC08pHt3HMorXOa2WUjSlRr108zODuXTCc27Gc6WXYqrVjp5+JItKV0um9KX61CP9xunqwuhf/5
knaZN6DGatTfzCCSPu2Wl3dmrR1D9yVeeCjSWRrMn3dHFAAn3zULtsvhp/NyoGoueo4/lbojTYa1
sHuMravjZzxBsp2IbbFrJPTuTDqDC4KBJasYnTCgfUdHiHxvrNjsN4WXhwC5CK4dbAsc4RLhE72Z
5uUVzrK1bHA1j7WsnO8dvUA40coir5TVuGA99rL8cBO74gPONZgKjRPB0rq/9Yj80m8DW7iPfOCh
tGsYPTFjiEBVJeAEfF7xbGDLyqtu7iYNwUEOJFZk0d4klSCHp0CgQYm7WrMHHfKwbwCB2CKqKdc+
p2olAa4BCCyA5uHDtCPpPBzRXt1V+GWH1uLoDPuif+DBjWV9+hu+vahqvWyoti+vD1BrfQ/HLQtM
svju9nzmcbgOf8pXJtIj7dMPFI2jKjXMLXYYhShe7Df/5YzWLyvqoSF3aXIlvs2lr0eoSGj+pmSP
ec3ie79R8dOZy6HNcGaZwWFTgKZ/0PrCcTds88O34iVkdWhP0/RtoeibVHNPEMOIPhJvWFTaHL2/
0bEzEwpmmKnvYXqOtAkR9XwaOTLRQieeniuZUDPlx08WkCu53ACnbef13Qixg45G5BSHojvdSM2d
gcKv2enOwK+Y3gMlh8x/2ToSWnCN4myxgqb1fAQnO/yx3KGKSqBw0OrDLCFf/4+z46YM4gS1C5FZ
aYABLgfkKfi78cLGmJxCYPx6Et82l2VUX1DoMHr2eJxJqQFu00VWhnOWTuBy1W2pSLjZSYcbK++X
n2X0ZdU5YihL00JdKAa7JS7RP8WR7mV89uJD/wngtZw9gvlfvPL6TvI2t7vfFUJ14NR+xi0Mk7o3
5Th4cS+gmylzETYUTSRwqhdZt+Hpdw/pIupbP9ceyk3kmYxKQYFSthC6QGYyQFxZGnz/joaNiKMX
l5ZY1rDNNpfcsepGlNYUxpdGwf9DKX6UyEk4MHHG8qqFkGBn6Su+ywH17w2NkmiijQ5VaEdFvjXM
IJuTm61gVn8pAVxwzA5QvQ8LkUE4o3cDQ61BjvdEg0z6dVjWgrllWZ2KQqMe95vDgO+EHStUSiUq
4sTkiCELMNAPyQBHsL0NhSzj4it5ZJqrxgJwD2EDrqexAZFGqx3a5R9NuuEom5W84HQy4EgsGeuO
JBYEtQYFqY/f1c156Bi/9ZnN/qXME7k1C48ecxGC7dWw94U7al3gjdaW4f9lUAjsbS3c/xUTWtHx
NhGAXbic/SPmEeb8REWk+XHC60C4yWFE0nlzIahBs3OG2DhfyPcltEnM8PlAgk4A6f7oqvSc67Ha
R7qy91JZR3qtFgGlz79uQ5AA56gXg68YBmFpBvwQSPrf4b4xnhpaR3K8C8C2xYO+e1LoNhzxsBQu
RazxnICFH5gS5k8w2ikv10SLPVcGuCoWjKczLTMxDq5QwZbPrKOldZURoh2FiGFaTiPJJFX/E65x
Dt7lUSunA0p/pqT4SA41YvgeOfBVKcwgcft2TQZsPmp4llZrNG5jRuevj9vk2mYbp9tMNYuM/Xxy
GxnKGy3Vsm5FVs+pbFo3BoRXbt5pcaGSOnUCeB0NGQqILEPTc4eeg31ExRZatXezWwnwbOUG7wKG
eV6EdnsUOw1DAbSEz+pDkLTBVqkRx3AO/CQCEvscDHmvckCn+YxPmKwT7z/IXdfNayxm3s0lNXwi
FWXqEIJGEh4OXky4O/vFMaBMA/jOJXPGGvMz4S/JTXQzI3F+bQfKOPm82bLWBtQjhISazcMDrfzJ
9WEQbVicSbO1FDlFzKYvWxJ1IpJ01DO113kFskHZdqyw37PeZSexAjpuimfMdMVPSsj9PedhQL0p
LYTMa56+7iOUQDTSFv+VpFh7oIg50AKATs2XVC/ZioFjZROOh21r6lJrZQ4sHBsZrSVMX7OEmLoq
0nKNVxrJ9NL8kCMoyDZ+bizqMb5BMlYSKu/txME/PlYDyvUX9ZsXOjimlUk35zsfvcOL6NtR/rF3
W7Na11KEORShwT6p/HJOWTmwI4kiTRA5mo9lRGQqFMXqyCQ0mFxjuHX1XPNpiEZdCywLgX4L4j0x
eSuZgr86r30Yf3WjkB088kyXuHKUfirXHjPFOUwARcwHiSP5rOaWWy7zK/8he6CJIlOcJfWT3Dj6
VJ3h9ktYwyZRBE7BwpRX7qhLP3TDPKYIk0QlKBjpyaLoyeD+KEiRUOvJztRX+dj4Lr36DzRWjP2w
FziM+mbwpG92WYEKk8n9PEPehjp+neRrSO02/1lUr2AD0ZsA6b74DGg5ydUvCQWP0UUPcjw6+akU
XhAqHS1U7wOPmylc8cmzjarIm82DPRrZr9PBACZ4FCR/6x7JWRrCCjsX7eNdQxTwvtvQDWxpMXSF
+dJuxNZwWTQtMku5PXGKuUJ/PTtUs9+kSLW65nK8op9E4EDCUxDyWzoY/UmUHZ3LBZJ/IsuuQ2mp
Azed6WHJLOJGT8fEgVnPc4aH1uWk1jsoPgaeBpCclBctRwJDub4LulQ1CRDYugqQEgHTfkB+mEwy
BXHRXro+nY1qo8cvrV3tDIYod/mNNBQIG0n2hRYqbZQPbBvgXeNnScorH7vGduOVqf/sif3lCvbT
KMInQLeC9NtTkV+L3p5Wd2FXqybuJJEgvGu64/ub9jwc0An3Prx57gS+wM36XdwBRQFAw5roNnIP
j3d9/mowLFE1Jxw1R40VfX/QMWeUzmV41z6ioCg9FZF4j0QEFKtsq8EbsX2Fu2+8+zE94wGnsyNW
z4Oh+BSzwJvq4foJoorMi0DC1X/FvwR+IxyJ43y7YZQnpM9KxOSopwcPJWgMLmVZXJzKEhW4XW38
PnTRgetyD2tN1akAYQEJIMTqfCh/K6fxPwkxdTRRX1E3F9ja06Ip/4BVxd1Vs7Or3Ftodu04bJiH
d8H7p/ZS1s3EeVvL7K7oOj6vzJoC/Ua4yS++yVstAgb5Yvc5BFPNniW+nNwtcr8Q1oYgCPVSo8cO
4zkiK7vLB+EqR/fhkuL+aFrxW4S2Jtz62/5EvdbiUB5rYx+lMS78DbugbnEBFftAmrHK1bDK7oK6
KYOVNG9EWUoK0BSQczkOiSV6fl74gqp6j6QNlwT8KiJ+PjhpwAXediNICqoJUwvUc50d0KrHJrd7
aLCG4RrtnKHyQ+nxA1nB1JEFyznIokH3G8TgFbBzOpKhD/qsyAzoe7qHfjx7YT249l21ptkRA5eD
ykvSP5B9LFt8TcuUOYk4Ck6WhvTvFRT/WS2e+kJ0JzHzNs+4+XgKl8kzhbv6y0STL5YLvkcLl8q1
glHW/xQdpGk8ynjnpy6N2pjEGr1wOQX/hzqkO2SyhyXQrsG/9pCxwcBp3/jzEISO8jBShuT9MNrH
t+NFKEy+84gAAvSPxbANg+5i4oKaKZov6IPkTz1M7uLWpgqnK5ru6UCkorhB7XNIlN5rphABYN0d
6Fxhgn+IsJYKbls6FlCuVLMrR1pa/nqovycs1TN4xhQQO76R5wEF8K6qX46Ttl1fqPxJn8SXs0Qs
/EAr0z8Rrp//DWDO5FOKCe3ycYz/cWO+wgf4QSGKvthPKLgBw/RbP0koxjDVzaIKniBGjhLDaJJW
rJ9iik1T2azxyP69KCfEdKzWKskjrtdxWn19Z5YcCd54fJPSusOIJ8H1sK7iQMx1C7udHb+ZQqyx
d8PLDmvzd7X4XxUX8/9ghpKXOIgzysYV1oEJcvqlDQGinT2YQV2FLx+O8nSvNfcusP54+0NLNpw1
4WQ2aX/CjWTqRe1eTFEubKOWlB59bFLKVplvo8bwBPMTY9MeXeB2T40PCn7Q/6VmUrLzQ7ofiMcC
j1YqCV10GevSFpc05y3NaEf6B5ScD5kn67whHuiJtSjz7Q8Ip5ca19EEnmg6nHS0l7Ds9HkGQXmB
s7cWgRuyZLe5khCkVixQYFQimARC7/k7XHIMSnuKf+vSxlg4DK7PVTsNBf/Xb5yIXylFKVidh8oa
sIh9t/LFLFpxx8eTAAQeRjxrmFNRaVyAaZa6YlPX4oxO1L3XvDA13wF8zoo8M5iCAj2EpV6OmWs9
xKNERXp66Z1blwvRkrn2XsaJ3QsQfnMXuii/w3dJosT8GU+pjRPZlgT6aanpWh0JTowaitWHB5Gg
UOZdZ+2Na3c/PEVFhBnZWPxy+APuuWJB5r5RAEog0xC8v9vJItAW5EFWdW9TvZ5Tm+mxhpMDPKLn
/L22U3CkraZWAbwl/CFKecqyGW5E5FwJ0obn9SxuXXsyX3n3NBGWPdMtdHws4P2OQysoNdQ29WOK
6Fn8C5FLRJdU30unuYRmH5VZkkPtgw8YNoVrQdSqjLFUzeDin4y0pfkKFypyh8rrRBiOPIEshaOO
7sUz7PUszW3OU5x3Dq5pnbd3ZuPyvMrhE6d6TZPkJpKsLgX7CJRfNYY/ZNUgd9a75hjgYIX71PJe
ZTsBzt30fID2fQJLfwKjxBfe48ZvDoexUDf4jNUV6P7yh84fd5eCSEIsYkCCkCFU/uHBpQjoUbBs
3w4Ns7o75Of8TM/oDW1eXn7mPB62g30j6JLkJxlip4WB6pwFPDBhfoiBWww5AzhXyel09blcz6XE
YJi5XtJkDSOTRGoKu/+54kXJZ2H5xSCI8/CT0Vg9I1OYyUzkLi+CaWX7gtYrNzHXV8KQSnak5zV/
8ZXO+tYNcP0xgvolnkJsM48Az45TpBhEWs+q/KXfaZyBmLq4X/VIYy5TJCROIx5H1AjEGEC8lkfw
1OnkWHVhDUA/QXMiAxhLZPI1zADQ9CTffALP4rFbBuNe++RtnUkOjnqA38mBdC/Csgxxbo0EArIs
fSV55+6a41SQTLkiFPw9DzGtHniBnMxjua7FJmeovWSaRsVGqrr4ntP9eBluEjjBlR75A2y3t6rw
X/MD5OgQ7qxnkukhhjGYfKXxsySVqXb0EHtJzaV5v64NM9W7sJVew2h7LLQV7VR+D79NYpj6+dyj
VLWp1iRDo4P9hdl6AO/wsu3HevTaCNsKcUIHQ+izFe3+ECyu3vw0KfzXXhvfLA4tGFGmlyn8MQvg
zmMHPYMggaZPGP1zbdmkEaxG6puar1gMlZ26DuCZk6i28KKs1A0ifA3ZrhT37TqwAaLRLp3DZ9l0
pCrs0LFh1qQFzIBIpv4ILPz930sKUoN8HbumGRZj510kr3pIloclGLHbC1LxztuAIPlB3GhVYP2G
sA5NEl+j1I9Xkcjl7zDQAoa/TWk/TvXytlNPkoeOqay3z1iP30OCR0G3Ab56KmN8FmdGinXGmPgC
rDQu21LlplMFKMIE3y7RDFWLoN/ZA6VsDo+t7f1JzUu7leriLEpMcAT0GJUW4zal6QWBIGq+QNSw
9Hqt8eX2icmPlTpxISxmdYWU/sPkFYfrb3j5UYJgDrMT+ouTCY/vQhMDRF/1kd/zu1LFX845qyo3
VqYaH+W8MUKowoJRJqoytN5Juuy0XKWPYHXoP3344h6/Ff7nfP+Duzq/MujEocWp81K9DTpIuIDt
lAjVUOJJXBeUE6x+z+he92xeHlI4MtSc3OmGgJcpdhAXIVTyICxg1QLNg4n7CKrMbc7f1T8H2FgA
mx/DOaMWH5sKPR69R4n6EGJaAb0SLexsGIctNpfEhr8DMyPd7ACit5NSI0yvtyHHmCof327E52Iw
ZDY+G5KLaAvpwHRYISQ0EOxlU1JCE03bI56bNgoeeSA2dK1aCuIxhmCEZQPVn15/WxHb6MF+eF5A
wa+hiDQA2gaGyMID2hceSqWabAy3w+3jSmpRRa/UDHPm9/rLkvTL3O2nX2tB2Gr8QdSCZRBWJvF4
qPlLWLeAAmnwZYyCo8yHGHXIqI33CxfW5gCACdr8++lOwpjI1qVA58359eNr+/3iaf7xWkOvi9Z9
EsZi3CSKgGBq8l7k2Mqmt9/pMIlz34Q5AKlbEpr4Hin+hl7efN1uGXvSTNq/r7G2EhnxqBFn7u6l
OUeNrZwI6WBecg9B9QfcDAnfU6Ta5EKUH4lQ8EcRzliblrnvkWC9egTOSL7ZVj23L2WdHTlP13BS
cz0kD2fat6ThZ0nXkp0B+Ynrtlyvfu5qbbKS5cuv+YNPlL7D7mTRpzwqU2SGNQk9r2jjq72rmZT8
9NA4skCdXQ0gEJkIyas7nhewWaOh4gHpOiS4esoTMk4+ZlV9xkgaUnXVZNZc+TXiXBfj6ooFIDHJ
SK/pc2vUV3y4z8FQNBvR8gEJkaKh3Lhwss/Q077nCBzlHqFsfV0BADFCK/yrpvQwfm6Z9xdMrVdb
W1yVuQ9GvCJDDOdJiTh61POFRh/b3NHWH+oxXyMqybXJRgcygwUNnM/hctK2w9wPnnHAuPKmrZ4p
dCNF1XKxYX/0TbtqKWsdO8Zht0b/7wSvkNjjxJAUq1IHoNWRA+0/tNp9jMNUZ/rvtusn1oUwD+1d
w8H+DBN0c5E+MBb8NDduyVp09Vfm85OZWWo+cyXRjOmHuZHtIAjdsZFLoZ2OguzfqQHI9+av6S/4
FgI940uQ4V6lVmfwN0ALSBmhzy3+o6LnWoc/FmbXW08CClPs4NGwUgATQ8njtpZVgvJuHBGKYCOC
o6snm1izNhw8UPVZC/yHCmLOd+qVHxCw11TygfAF1hbDZhusX9M/uet/MEtf5xD8UH3CBXdrqNQc
xiLyAizX2XLClsNsZay2jbkVieEGoXEn5O9a3AWu4eUPuHGar5W/WBOvzsSESya6N0QzbWMz/rLu
n1gpf/jLGBMtJ4YvNh5gb2ZCsgcpDJvaOfI9oImo5fiGMmEoQlaCn+lsOEWxdb2ZIlvkgfENSSlE
lBxD/odGHofxeeYJuUrgBS+AVb+oatGekbI4sMhp7xfxytG0jmWs2RJ3Ck3XFwJOutkk6KE6dvm6
Jl7JbFYqVTB6gRQn8YnZDMHl02ffD25xavjgv5ppMtkYTSuxVo8CJIRV73feEJSmkYucOsgFa/oT
01WY9AErSa7PpEXOWmQ+4hM1y5SaLGZ7uKvQOW2MBXvFnYTRRqGKfTy7zcBed23h+NuSsgMZbP9v
FsEJNEE96AvqDKwHF7rfQIHBv9a6OrIapYrNbGgyHeLWH8eHXl0in9pPcqKeSmqB1OKSfd9kkCr1
UJ/ArzGS67lInzlEDsWBqRELSaXUPO2dY0jKMHhFwM08dBJ0dcz46OJxFdOXfeMXPf6i6RLQRuJc
TjpwJMaXF3vh3HFhaNkK2iuRbb0Y5dgZd26qqLxmhAzQ/hFRR8futjUGA0Vy4bGCRkaMPtaXr7hO
q7h5bRD3P0cRVKLK4FvZYpLaf/8DSNcANiofEGBQFML2ROwxbZPonlO3trf3I1jCqwJZ6TmCrYl8
vzdpsQ8Q9NJqL3P1dKv/5/fO0QupIXdMXBcu3pR5J/JZfPx5qqj9kL+fhZw0D3H5t1nhBi+hfqVT
YhccBqB4MQl0oKP+8sQhxm29VNBnFfMYV18zD98KJ1B6xS69CWyofcnS5eq4WXsJgteOB3fQxGAj
gM6uvu9xc+bWY6Hfpa1P0E8Kr4T5orFLWQkY/ioenmP/RvisYUSV+Vg/daqsjwn0lNsnYXDcByis
enDX6tqVYGgNTPRIM4pBfmIo6JiJxSTvJRhk5yaj/jdtszFfhJSLWqpuIrNM7AmL8CKmJyzq24yP
pnOlxlX3gtMaGyu0xrlR1+Btyqilk9RUfbo1qjcNwkr0CxgvlevBmro656SCvCcui1unUBlakbN2
kxgaYD63kzBIbe3wkqtGQKFvNFejdZ6adrC7KVZdM6qfRCWPlspxRsl8VVYkNQdyYhPa5m+KXfBQ
PB0vrhukoVWZ0DK10tEOjHNp8eQxU1CBLb8EvTpYvUnI/5BIgGwMpPa99+CIrW3xbt1NBUTZqH8J
yV0tL6P4bh5/ogrkcHy1bVue8sq70Q0vvkQNdku2LTrqJPX8A8Bpz8nigISLPtXsMVYxXib/pZMB
9/7hpcGqFBo3imO/AampV6MRkooqiMPrI+9hzZOM1oSHsI0+kv9+mvQl1uQHFNWh1cjwZ7MTHxks
KlF8xFhB73N+C9XlwjSzyR4abb6Q9xPt8ZGxnJTRurYtseqWMwY7ZwBbT7fZIKFGQ37L33v1IReg
KjLf/ng3AGx1YazjjV303GCkV+rTo/CRPamkA7goZhAWgxdZQnOfyDwMPmkblvhQ7OXJNRVO1705
nCNgrtr0oxz5Wi2utmHsLMJK+Fu+uLPi8dZOMGd4S90WrHyOWZLwtuscF7ERdPc4e4bus3JTznyw
iieGcpDTRsIRaD7iUSwTZ77gqRgk0VlJXOH8W83+aKUvyAswV/wFHEMgJYl73xq4h27U/LivJrXy
9RVPmIH+cHHiJxmD84cqV3+wGUiH3a83HsR7aSyQOw6+G9/PHKGXFoTqSsGJC3jxzs1NS4+SOtwb
0RTBTqQ6rQgERsGaNpAHSS/RoJnti+wDGt0rJEXcf4l/2eH3WNTLzo2uN6+zWWHYunAtpkOS/NpP
lTEUybKg4Ys0Mgk0WgWqNWpCpdZg/FyGryClTCJi62cqdLXtbJ4QdxI2cXa0akCkPnLsixtINMgq
C5YPKYoTDZxraVTQwSHMsF0gg5OmgINeIWArUTJFk9Lvp0NtiJIngpPqks1HrMgaUW9xkrMCcVzn
lOcVHDr1iz9875pH34dW99bm2BFK1w8y8hiPCCFhbY6c29VP4RM8v+Vgc9KPmzk0XqbO/QOlRby+
+t4kNPtMeZa342GhP0aOApJI1+ynSF7BwOkW1cHB5gJbxXvIBnRyiiWpgGw/oksHe60AvRjXK752
6FeYowS5qv/5EBeWrdMo7iJ5DZhrTVmzgh0xiMPC59o8K+xyphPQixwhyN14yvATtCvcl33TY2rl
XIqZrNhla/wOP72Hj6laMtAiFxD87zZhR2cZoud76JRxOn4JnH7Ym57XpbXsrOxAkHC2z2Tki5vO
KsMSlpXIGnGjaUflPrjvFbGhal8afxoqsp+mE+8+/Lkm+5+fQrMshStr3XVNqCEdgRsKdy18XMn2
Ph5GquUMXxn2bBr8AnyjHHm3LVcCLI/zGD6liVMkHv0eq3yQHTxPTtZRw9AdjyUhXMb8tInG5E6D
UztXtya/6YXk0EZEBJPB4M0na7GTEem/tTVWz1tG4X1m1w6M5EC9RqA56SS1zgoGQdfFtDhHRV9p
PFCuJwWr4L1vor8Pt8EVYqdnT0fYNwHA0pBhtN2Nr/yPR6uVuHSqTwjA1ED93hbDpGSYAKNVRVwV
A7+Rqm1ix6Gf9i2+/Ou0N2L56Z4StsydB9SwVBFyvWY+BbJFGGP0hC2woyYYMZhBEVXAR/kNNkPS
c7MRFPXyXpJFHcXiVf3I7oltBzZVqrjuohk/ONeJzHBB8jFUwZyYtyMPYONyPjX+2wYviFjgJLYM
I6Q40VzJOlQn3TLL/jG+RHPiFq1EIR553N+vK91Tj8xf+u7wbzUOlAM5ZAVJCDfMalsDtZV434+n
DGohks47XIv18G3g2IEZvFL42Mmra0DReXU4qIDmtaqkCFsw3pkcEtHFfeCaNxVSGs51ywjc6rWa
g4xq6xsjZJc3eNnTH9B5cyZfHRZJ82QQ7vvV10TH0XhIaQTVwrwM7PRixZHzD9+OKaneeKFfeP46
X59WWv7zaRO2Wh2F3UGYa/A2v6SHbt3X+5OCkAGJqk21FHqwa08R1MjFle0AfP1PbgLARNus2zUO
g2Cdu5kZc8cCTnPBCtM//sV7vyEdAPlQeDB0eTeVO8C4asyw1OYVhIOQAZagrk5hNRXHEWlxsPCe
QFA5+UDFsRlS/gVDnHkI0qbIk69lGkBY/gHNL5BWk0jD2x2G/kN+8WXOstj2lbd9FC9kImdZMqH/
ROHTZ9HTxE2hxQVRmmnJ4Wki4gzBt46wqIKfyj/qGOXvX/1iWvR6V0uJp0x/3SdHUA/h3yz6vCo6
gSJNN7sJfrgPEKXLnk/c6d+/hhqrvaWxQKc7Z5Ica7pGePb1nMuJwfXpfiCTrX5jpgoM0R61EeCg
0aQ4X2sTM+diQmuxC/atbpcqfq6CUdjowBgUagUwjg9KOjSezz8dwlz8fC0n7qGdHm/YezTAoa3C
1onw6Abq8bwxmJeOgt2s31UUHsI7PE2iKVkhtEBHYrH3AKCzcYJxnnrB/zzCn603Sl0XYbwFXu9q
t9Ddmdu1Ks4p1XYq4EEURyMZNr3vmlPGdA32HxtECvIKQgf5vFx/uyWLLtFYjtE5g0f50PE8L8sV
IJAvSgHdaz+6ZrIthWBSEdNhzm+ycvuBEze6QnW4YKtBJMBVV4FXkNXpgHRgdSbHTHVDTKGnkjQj
ZZnXMXMJLQ3dHyTezPM/uRBf9yTboJyGAUz/fL0Ruw5ma+rQPGJPTY6qrLVqCYei1TP2Y7nfhOGg
SOFQSn2Pht4ShIgJZQKryNA09BUbIY6tYG8rP6bOQy2Exx4zJFAIkefyZ3rcniGgx3nlQnxG3B/l
LYDU+FN7FRLQ10KPjw+Qp/vn5spUnWOwt3M1WRO8PUyWWVzVCVSQEOH4gEd+yLKz1bFKZYfx3huG
X589FvJNQJ/hA306ReHeD/dpzeuSsHeTF7bEO0HStw93FXwQ3TezAKVY/82Cy5WraqjKlQBtgp77
w7IqRZHMXAinniuZqoFk2xSk0L8tbNMMml7nIVkkV95jqas4gJFgUPgUzbW5wirxwVXaeqa/SQFN
TFxrpkmeMin01L2JbGjaxV7V4atPEb7NL5jd6aYsJzavfWAaFb81IehDYvblqyHK0u9IJAY62vc7
ehCaa12JPKdSWI+R84LxtluMmqiPt0Y4WZo8ni6opxjwYGf3f5d7qN9d+ZyNfz3YpBiMiew4/y9b
YAMNi6dbZuDmDbp2ST/xIqBH01FXxtwa+smD9+7lHnPWMLgUlRk4ro3Vu2BuMQJHOrQGOg/xLjAF
+Zk6chX1zaiQdnMwZueuWCaFLcuVJ3viWpDXHAbyd5BQTvvj+l31ySCyUt+MOLMSvDQYJWUQV0VU
ALiRYn2C/Gi31n/rbQhjVTey0cbxajPug6TxyhYonKHlc18D0dPEmcWx+gDfcoxUxPjRK2ULZ6Bp
fhay/4uD4diAzkQM/0hgcZL1TerLeUtmHWVAAC3CI4gD7Xlm9n7AtABoht5OekfTouutacm3VoL8
nnpCmShN6cxj/zn8c8HiEKJ9gm9vF9azK0kO8Xw797uawhbddk9zrDpqEOkD+kA6Dm8UbNfx/mgp
wmAJuyp2qq/uMSZaXeRc9l5mBKxVHND6ghiuqwPCq8iS8KP/L1SAHBvd6/wKW/kIrn7Bj9O1mUuB
9zMQaDFQfc3jj+XHlL+ums5tao0Ee0KDQs6onVu2W5XVGvf3zjBNFD3B4mqYswHqfsDSOYuVoUJX
HwHa+UanBco9RI8E2QnoEbSzd+vHHTuc6zATMgNyL1IfynePcsiN93gNzTJ7vmCqC7qMJ2t99N+I
WvlMp/89T9mahLe/bxCHZTG40WrhLe3LPvnnprqZG7hFe8SSM9X9C2Av27i+pFi2zixWvUaryB6x
lwKWx1FINREZ87eJ9Uc8eFGDWg5RrgSLIhyXxoMh3sv3ZsfbNIzGXzAmlVvTgl6UD1XoMQl3Mqle
EGu7scKQ5a5x5T4RXwvmoxu2oVgob96mAMGbi0EITfzDefHX/YR8N5FVgRpLALLS9b6Zxmc0ULwk
7FOamHjN87g6arCkUAdWNhJn5O/ThNGVe9dcXY1yyo8pQfUefM4xCmFy6Kyrp8JajWd+0loOnYcD
W96NAzEhPxjS5lnU1R2OaaDE9sMwsS+73UpIaJBwuLnNzw5v0TIRnw2DoWKy2fnO96ehmEHTqQxx
YK9PXhTCqHeQJOqEUOFxihnU0pLS2XG1xHc9RsaRPODm05rPchx2J7T3gZT4Le8PVI22xHZ2xZop
zeRSXsCV892FojbCY1YSOxGhb1H3ODZjE2VxRhqmLoahxMEWL6DLQjWyEyjso62hsFnXUw9c7wWZ
r4IURBlz9SqNI5/D9LZo0l9Xn9ESZGeIUb2WhJNdecgCKaNL0s+sWO5y9ptTovyV8t4kRz6AzELj
kUjEAWL7RulQc9lKMlHf0BuGJlsyIgcOP8UZKTBCCc11vz4SJuKyZ5G0UyhNXkk6c7DX6Uk3dk5N
tvfuGsfhLQzmWG9jwnPI6XZGG36e/Y5b+T+rfxXTxJqrty3wGMqGJmV1VppAgd4lZpXHDGjRFVzJ
v/jSqqNpFsTIZimee/0RRQCn5TPTVmZIS9RKI3c10f5/1PepIjuci+QxmqUESx1G4Q3X0SF+gv2v
sQkxtFlKlvf5XMPgeKdVRgLQ9yOyqbUg4At6QOlpmE/3Lu7e+iadZOGZ/qrtrmEz98ZdSXm1InqB
0fM4itbWs7mko4Kc+06AJxP1hq4xUPwhQPcuV/IV/CYmPn/rDcxya179Srr6ZykrraPM3SzvTDwe
6NkacP6Xojy9q5ZNWeXV1fWna96WsiQbTySHPqpyFYOHewc5CQNSI60sLzgp9YLqwbozeB0l8I9i
CmsSfaiZ68DJsUwbTsIwREt/8HHaU4JxjMjO/dG6JVM+vrmckqJuIERC6RFwm533ab0GGtRg0fV5
cK6BvBZkNxYDldhXUGLSfkpmBBGMHlem86afeSdo2Qs7m7c3A3l6lADE3vLbhS421xEZuY5z9zAg
Jexu3o6+C2+E8qc4l1pZ9qs/O/7kpXOyJ9X7KzNixR6FfxRlwmVTTws94nx8wnmOy93yjkC0nfEQ
AIix3n9YzrChwfheyp5q1khq0FSn0ZKUV9Ni8elP2EIJ2SVL+AV647d+vSd+c0MW9SLEAbYIfp8V
u63/vpc2agBgxu6b5592v47y0dlNWXDGi8we0bef5NHEKSS2B90rg1m50235+/Md4UztcA+l+JpJ
c1pM56TIBOsM3uViyhZuDhQNijsStVhubNNIjJSSMBDIsmRsulZ/WAWZ+2vGei4yXY1AYDNt6dop
b43mU8EVRvpl2qp0Kq6TOB016R5Ao5yXZycInbHXjDbM1vkYXWO2A8Oyj34AQ1vy8hlP3K/1keJs
7wfnHnlAsNHcQzT3GxfeJE9diS1DdhVUzJ/ArZouieaPCOKSLs5iXk/c+ZfGUn2Ym0sOlRZo8VhC
Ltzxbyxeo+g7b845sxD2Dy6OpDuzUm+ODsCwO5Zh+x5my6LMYobaYDYDbIyeUXfQJn+IeCZBDjxC
JP3rkVFlzekeauDzfGF+SM5WZsfdae2BhcwuvMFc6yt/yd/WLUB+p6/pcEQF+Nqz6MuZj9Tnq5Vc
YWRMqF0V1H/9LkFLMEH5naBaiZolTzaYl3VDGJ05EOpvT+XaeBXALUJq2ebUpa7zuxGy8xsm5/fk
jOoRPAvRCAcEkzYcXbHyCgJ3gJF3Qk3zwAUYFUFeFofAVxZB3fBcLbVxus1pKIAAY9NvVbPuC0zz
DsjSrQEtumSwVp9YNKA+SbsRjdgpRKFeZiIgnPmrYPK65weS56w6mwyZIH4evnAH8ENrcfjO5I0p
MW5npzqlYVozalm8CbwndIPwRSjChN/pYG0l8YgqGGBqN8re/RPxNkKAGkgqDytZ0aAlJaZ4gsta
zBv1U4C/uCDdiFszMqaO1k2UrG3IhAJiGlFXnHRDmpDV2ZHWWKxva/4SVQK6+fY8RK7YTp66HO6m
onM22/yFzYoi0wKfU/d20+AqBblOwum1eo/zb5ULF9YNdg7d1nvKsThR0QEMg9n6+g2vAqiewW6V
uXND3cJmyObbjfKroIEn+JwKse/iNsyL69Mkt4BusRz+kstsv9PkKDi3p8V4Bs3Z0/8x/Gg+va72
yethQ036qy1QEvqnSOpJVLeGbMsbmXytllefDZX2VU89Cn4N8RbQGmVCXCyBNOQ0eP5xyKkjXfu2
Q4NDfgxHw08h84WVWsMTMmfS+BnPcqGP63L2jbY8iTT226if/QUqvcb53ahjb9H1UwYm2V3O+BHt
Yf4QnGyFrb3fbX26LRdMvl87goMFFAcDezFzYhTZRzUj2I2w7VnZPTp8ZmUKpO2DHhecMy2SJa7D
58kwlJ500pM6qkxh/6djwdRSKefkfUlKS8COxix+5+Bwgo5El1/WwE19gSiKbELLjKwVmE68iENd
Y5AMciioo9SZk2mLYokjIcd03XX+aEj8I6SoWxuxU33LcsK+xy5i9qbdudc0QeSFEmqP04E/4+Ht
FrUs5uMozAgcyeVrkmYJxfA83NtSYRptgLQBB0bVJMXHGYCJgzTf2z1Wmhao+l97hZ+4NG92vxzm
zTp85ogPCSDM8fEUnpq1Nm/jkob+o8AI6WqOuZrIPu2rkHQF9UnXXVQClyFNNOnfE0+mw5//456G
l35N+Jidq5idR9GyPUVpgsxu8tlMdzC/7rmryZW5UJc9IXNrlpCyZvNux2IAFJiE6Z3c55/5/HRX
xcZ3kiAQvfxqXlb58+oYkFNdgWZ+5QZ5xK3g5rfpTAS/37Tdaju9QEf9nkHGxU9P7yORtS5BH/hh
cb3Rq7JIFM/nJK5wTFgO1dXZyrQL1XsshE/AWNy8S4Y+IbKjZTq4IlYDhtTm0Us1GAu5SEKQ8Fr7
nvTA81YYXa7tWnQAMc+Sotk1g6L7WqqosohF9fa/v4OdF7QmyR8hTfNMC/9+oCM8bNsPi1fOZJe1
yk6nF3iBed8UXHEQtiG6GdXFOFadksApfkfOkPSU0iCpAqCDgvjU4OUooseq3Z/m06JpEF+9SWCB
KoL7HczvVNLVKSpM5OuB2vr3nQVVa3zbBDTilTMO6GadoKh2Jm3CS8zp1KDIJ8TZxkbyi39rsi8Y
I+InbBJRKgf2erbBOdFLhc8USWw0sD1J/r+XhC7XDCvmEfO8CRP9Q/q50lui21C9yeP6SoUCV4Ft
CkEiEeOPIcfH7JhMooStiWKcOyH2DJTFnsJRYQcP0DOlTfCQvmZR0ZqI0332RmVZ4W0WWOPaxlnp
8mvDTpQ4EjSwOQHE7A5itjqCCT7UK6F0We52Gg+acR3CWMqGR2zkydO+gIbNPiVc5SI/gJ9E6VXH
VAczOd08687Lt3wPgTBIBahNoWoNnqWOh6plj7SubCbBXjSK77huNsm5XQ2DZTY4V8FCGMmp1OzY
i7UMiBRhvT9Jpn/la25oGOrSVqAWju2747Ql47+/HkljILWtM46m1I708V+Ab3BjV1JWJSDzOnUS
MThhqLeW955srhKTFSMJ0Kz6OAtUVMUwNkASYDacKFju9xtW9/j8PYFYIirxIxn7zpn1sfPmtXKL
+bUVkrqBp/eWRRikXf7Z+xYYlBUFep5hWon+p4MEIK+A3e5R5V25FuGDOB16aPrb2i7jzgT6q/r4
tyjmHaMGhAVLHuCfV0JMc2u+CkQ64rRRMpNYT9Ab5BGVA75x+C5YER/R7gUEQlTAtaJ2pxGoGJuc
OqiCJzRZxmveOz5JH4/wgbXqdFNU8q7puIlo3ehFmO3y1LVUueYtOYKHBCT0ihsK2U8RnjL4CZtE
pLrAQnXUhpDkAoiTMHLCJdML7Z/2JEMsYHlMTdWuMXQgaa16eLG93WWlSstT2hZl1ALjyno4v4ig
2fQsDhB+9RstLzfdZ1vWm5OMza4V9tN8+pZB6RJW3XWSHJJYkwaTOwgREi7oSgyA40SllTSmfPmQ
kSJJoSaC/WEI/xN/59vRPPe5zjRTzd9KcnXL6UD/4ASMo/8cScO5uy+5hwFh5sGeR/70HF2qUh5f
aT5hvAqG3BQjzoYgmSNCqvJbDrOflsn48oNguFVn9IH5PcowxT/1Vl1h3sYE6zWeAfMAlw7B368F
0B+aQ9knxjnsWEUrKEIEMR8mX5TaaIiIkek7va8we1AsTftBfluV2PHUdf6ThqPdMaUgchf8pyLS
5ffjfqLuxWk4JWaOfrSs4E78HZ8ejeVEgZL1sITSUnZbktxV0Nuv2OvSMwBW8JUhtFLSmOTuOyh1
b4n9xN/hs2XIxSubh/+8A7YKHKAawPs7nCmpAIQP08nRAFPlUm2dbhAjHcU7ttVWomAAAvHO5Nri
9acXiFwiiaGCs6C8xECJEzj1lBBqdR9FPvp2vlnJVn6k6Xbw4vuzUH+bKxe8C6ZfXvZ6oTDzLYL8
fz/k0J49WlClmz6R+vuHZBXtxr3NHJdf7OFzL6PmPYpo29Lz0fEu1X6LeJEkfxyZYlAg1BDNqLHy
0T+rgGBjI80xE3HN+v/DiJaYPMlqmHDCDl6otxE2xvb10XKu0rIm+UgSRzxRM6qO8SCe2TdNCEAC
+JOPSGZW0iHObLgFWz9ggJxZn19ijLMP821Us5Jl1Up2v7L2nHyNpWUNxqdUnZGpL1OH5RuAnHWk
nU1XBODZLQKMlGgFkY7Jha99QEHwzOTwQkFn3ZTWO+PXXHRXTipEd8kdaw8D7WVV7RLpoclLHEYH
C4SHVV9MeXHDqe3XmuGyGdlbYzdMXf01qT13azLGe60qzhPFMwLrBHGbW4a/d+2/jqcVs5qFlqSK
FEDDxsCYhcAY+FK9YMhMzRE4jVEGjbnwjLfpxKKZc5m9/mB+eJQC55fM1KGT5VYGkmSi5Th811P4
BOv5XgYcdubKZVng2iXwTi7YcGDeCgNnb7GPFnJ7k9AfjYrG7KnqC8b4WhyiAg618PiG3wlu73Q7
MmrE7R9/95pkh/bmUbk8RUQQ55gj73OXiGAh8SymWV15Y9Awc5pQUuUejNTdwiySu2Zd2Mkra+7y
D71GaZEO9g74Dzvg7p/qQBfOmYT0agZsv9Gnfd7DGM8xxTCwXQYWiGRDD135Pa3HT2LGyImzw7Dm
qsxM+v98gCxVx+ExxxYqI3RoXZmrTQ07jYyxFaEGTauUt2phUglOkOCqogROfP3ucGKxlIsSc1w4
K41/rmnSoZkK353FLYlhYTaYtwUGUISAm/z6E+WilufvgdSHKQHfeJCrH+5n88HRu/69foTCUnxF
Ct/qMuPi4nKWGJgPPlDuD/cnb0CI+0XysoRZ0JGAfdlep9/tqrGCq3Pf3ELLMCoU97OrZyBtc0fk
9dQqarcMipegPl3ihr+KfnRHq4bZFhy2lYdYMFb3DOFl+UgslGC0Q90R/FdnNWkQNPkE9keqYGBf
4IRBDBzW2kmzKg9EZIAWTzxdVLVtti4xhOHotluyuAOCEy8pRJK6dA2JMpHsxrfWMr3DA9e7mNaZ
j+pO/+HY5vTIWaAiKBRjKZ2Qt1oVWPWRMW9LfLPulIbDt4BTJQfsFGdDI2n0kBpHtbmt5HMG8yUU
6fHxX907E1MGtCRAsLZPSqDWkPp0FvGXdo/oV4uBlVPVVdCazldxQSnjdhFheB40YHGA5hw3xdZd
EBMunky9ENE8A2liBiXGj7fH4IooTsUElfr4ihFWHn3UFZtPG7dWivR/BvgiOjTG5ZhakwdBFHtn
bw5Uy2qf0YugQsqTE0mNl0Espxk2JjWwEImxOORLpjS73PrlI3Ng+3rBjxlnkpSYbEL8mvghVpKr
NJDXtayHYgsaPIJTUN+mfaCLGIRne6SiZFuHG7ByGKtCMu1v4+hlXwZz5y/qhAoIUfrYf7ki6u1V
UERTul3xLWj5Bj6pNsxuBYqH8T7kUFqpnMCzqeAW7kpvKTSmynt6UYBaIgdJaoZOk68dmcK/UO9G
NX6aJnYcCT5nZYxXpmQqsQ2ALCJLPTkmAXDeo4DvUvUpNiq9tVIDuVAmEZR315+Bpgq+toQlZp22
Yx80PuePsVtf2UXb2OvxSqE4JapH77ZTI262C9Up5XaMxEb4Jlz7mBQpcj9lsNDlPrA+TYnQlkLH
spdPAYfioxA8P6VkeiikVXqR3v+/CfKNUEHVTyG2vym9DaXv/1WUBKG4Tnfq+ufOC1DqDc9JbQNT
b6gYAGV9zx12dr+i5nWP6VPzdoWGYk59hDblpiCTa9nXR+Q5N/F4XGspt4tubEv8JnPJ+6pMbHfm
YuXDTPtVT3dhDFdX1e6DW8lDR7OstTGX6R6wvOWJkZ5isavCHCy1ylJZbZalT6Cr5pjMX7vdTT2N
1IYo91TyaG4VWZ57fYngjnBHqUdUr0wrxFQPRwIF2PF09HRiVwI5vk1SQzc0rkfDmV0tDfbF0t2s
6MXpCeEIlFKQJQABqoMXX0KpmaSruE3hYYN2fkDzb5qx0qFZPeaRuH9DALGSnvSaq8T2bNQo0m7g
NsJG7DKqEY/+yiiwXZ6gKE9/oIkhM+M5QiQcWPY9axwsro7utqz3qLkwaSiT1S19fZewe65LbfoB
QTuVfW76+nPVrcX3ccXDaCfaOiTblyZspzvSDMUMRGgU8Zws+LMnGvHe7A7E9Z2ImHgdxpWBgr8V
QgRXojqtA5SMdn9bjSwJeG3P+7GQM/nLjT48/lAosaNU4PB4rtw0AWzt8K26a5kaabym/MVLLMJw
pD7Jdrvk3SztM6m7J9V9DAW8QffRYelrbis82UERqkanyDBBoYoWKtfQVtEgcY364hB+S7VrI91X
AAEjvGz6j/yW/C63cj3FL+cHUbVnbAAKqIE4K/p7GzG8mYbq+OnYwoqjB55QfXfQOcPQ5+HXTUy9
VR4LXo8GfGSKBUE6BWtlEHuwoi/udDaTpINvXoChQ/13nTSvr11DMpiqjNzO+8vALjEOV5Rimf+5
00x8qy2JOsyEAV8yNosn3sBndU69ZA6E56Ehy3sZHA0lOAxxwYgFzehmkOpTraEcYJhespRKQpSw
rgtdUrDl3oq+PBPk7kYi77szV0yh1cz/RgkX5nv66kC8lGa9FRgc0DJ4OoUAFTMlsloqa3awMh/G
bditAKSwQ5+U/AHOJ1ELhmBf+YinJetLA4intZadS8PHGgPO4mPtO2DxKFvED09P5cEmjgoYvLEF
C5MlEbu8CLvd9OnxHuKFQ3AgfXTCyQ2K8Buz3kyafVRSqS7t25aw11Gjhvh5glrYeuf8udZI43er
OpQXvhc7btnrCOYxE1lCHOS2gEik3sdOY2uCd+CdYhkuAl2J1Bj2mNcjcs2GZiVZrhP0qpvD6nyq
oM7Ytt+E6A3glEpiAVzx4qP36eiE7Cq5IF9DSH7XBlBb7xTvSy7YJ9rA1sMLPd8fcwBm4NHPBB88
TlKf1oixuksH58NRcMUdxve6mwHpRe+aU4bzaBnkVFKhICCrEMu1tUcKOlgJVgRtrN9RCT2GcCPj
UgHRFXt6W1lTPwFVGsmIZJjtzzTTIQhgnduOuPmpkRsQWs+s5IYlcB55gYWo51iVRnoGhVdu9Ylt
PP746NcdTSJCAvQ8GDj+zeDf6R2ei6Eu5uKB5nLvrh798yngp8YclFbSq9R4CceSl/mZLf5jSMGo
8BdfYH7hQDhzXL8K+eT0RuE5N6SjhXOlts57QZBLEn5LMoNuQS/oyj3lNwsCiUE9fb7/eownPDJu
iOKudtGsoTJ4biu63/1mQFAJN1f79a863kA5aOS5iHdNbZLCFjxtt4DXJwEKTUi+M+nyRJndq8RQ
EUWU4glpSBXoVY3xIyAH5jVrkpboJmlrjZ6/tCrhzmkHWZFhnYXRtpvgsUgMIJMAE/hfY6RKKPWh
tJWvasr8eKBjvQ8xK2F3MrMPJrplnQS0/vK4aWzaBBzZDPCp95ASQC5jTDxqNli8M4E3OmjninXK
CzmDdO3+nsQHkSSTak2dXOU2Dbl0FfX00MLBe3b2e7YfMdfGFPl7A2Wj8Vqlxu6l/itKEygl2LMu
WUCOmP/PcDUkbC5E+CrpCA+L2y4sIvwPjmijBHhqo9uStFabU5ABeX5a6H0ET7hL4DK7WUSmWLOy
ldFFUCbW6zWnBKqof9lkMEI4xsTgCPZ3Sru71Ipf4f1NyVa8RPjG6AXyXQ0sOm09aZK6T/d/Nglf
WG5wP4j4xnyyPZWrsW9o+z8AFJGk5UAy26L4yEuLOLQZw01lAU6xBcEdBlQCKusdOlmMXq8INpSP
gyrXbsTsuBRN6W8wbAYm8sHX0QH+Nb30QP/DFCizPy07Qh/aBfVWhnpyscM//1oynWWVev65XJIM
ACpGB5IGDohxMALTrHVKzTN32hoZLtS7kYDqLgr88cqVNOAZsC8Gr9ZZiJpOqrAh0XfU8Uq7tww9
GLOOU0WuVLShrrTTUKE4D3DqpZhlSgtLvtejjGFSmASMPm+Hn5uPZ7X0UByH6zIqAXNe5NbYYIu1
TUEnmtXn8OVqHpBI18AnZKeeeiaBJRuErqSdMTTZTCSmBrKdb7bhlFb4j8GShXNMB3glx0M/F7ZM
rAIgazlYh1KGXnSISaWuxY7or7Q9nq++NXccEaLBZ5gl62pS4pxu6+FxksfWyjGIFntJKCl32bpj
XvIl56hUE8K3vBDHSxKZOOohqZJwwvAWWnuwvi7rtvCR4Cd52P7mfFhqrpL/I3Ua+uZV1yomoc4B
A1euy5CiMpNAG2Hd1niPCOLNEJcAejtc/5Y2lSRwSejFPN/pv3UBhxZskvkTKqpepz3kzYlAwMra
gb+rDujcHuukxpe1LxIGziotES25R8YQfr7ZGnLl6npnvbF14P0OX+7JW7aSPrkcmCKM7MqxJkhY
YBO9WbID6k/pTdn18aXFYdf/dz8CYaf0aT2XluoICft90K6M5gtrgTjw4KKjO4Lg5S/AmkvJJGxl
/LI/pGLzETfDhXemiYDBorBgUYtR5LxU2I1B+q5+54vt7H1+rz3rMlgtlIFQ5pR2ZEW3/dLzbHaV
ZCfJGmw9a/lHcjk2cM5BaJ79mDsM0v3gQCt9hX4wWkiMDz63dVlmw+LdvihZHGKNTX203vUWyYQW
aTN6b3t2fCVmM7+i5MoAH4h17kO8WsXS7odlsXt96kqepKLGJO2oWkk6K0pt0uJoI60k3o7nvWyH
YvPmACpCgqg6ge663x2EQM1I75kuX+0kHN/+UkAH5W2j/e0n9tCsL0e0f9yZXiVXf1Sgn5nv01fU
gwtD6bjXFvym34hGqq/WF2OM1UB558fj5wIigxb9IVSkSRRLUTiIAIQOmsbSpVBMdsuhsRoASfQn
++8YigVYca1sVtJpRA7AFr0k28qvzL3Jd421OLHU+jo6vL6x4/XQzjhmg635afNoJn1Tg5FUjYzr
zW0ElmwaQgQZG0nHLHW1v2EJbadhEYOIJi8eQqIh+gfmjzOTJginF6CqBe+iynZCA8AWLQWIdUpn
yYmxUUPwG4q9COl/E+K6imvCRC3U6ReN3tSN/Gk63gwgg11mWNn3OxuoVYp84xrusFNNS/RNx17/
1oKSTdItw8Gs+958oU+55ZSABgaJjFMorRs/ZVCUxSenSoE5nPTvSHsGjeHFvw0LZQ33BfPe9CGF
qqkDaCjjq9KC5QhEDtqb7Py6UTM2pIg729P4CMvLPvEIWAfkck7khtUviZI7mIDYDKGPEfZoWr5Z
LYlDSNtcj0LxBn9kC69fiYX2JCqVuGjzi6zPKkG89pJMjLZqycCFER8/Rs2mufFXTvk14o7ZOnU6
eYjATd7+i5cY2eHNftyWEHaP9j7lN9isKPjoNq9Xbet9XdfZSGNKI1/e8gfay0+sqSVR2nbUORUC
hURzavASk5RC7j9VQK8PLc/R+QPtRrX82LULMvWpDAc6pY0Wt+f/jWfWaGouXZdpUSOVH4Hwnuol
HtCoOMwMzGXTp2OQaw81cVKw6JlTvAhSN83ozHV2QBQ1ArljF09wc43ATcqbSC+j5ZFkobz/r3E5
uCd11eFk+znmUj9XwHUEeJm1u/OLJET/1hAbd7Zgr6q2Y2eODMg2xpbi56alRpsxFUvtQPJxxFPN
zEy45epfB86CptFOTX9iIl7mOR57uA864tuzAARaidXgx8JGptHaQVh2PHHX/SOdc6FdHkSa+nLP
j0mPu/+DVyG4+fvCVO2S4s9NRMLapQ6upvkwz0va1CCcPLxANgODBdYg1j5Lm8GGy4NCtf6W/PzJ
Pm6Qg7e1FgbevVJDFs/AOczcma4vkImqWSDz6WWcXbHC4emL5iuJjrEyuV/K7Bax9E53k0jx4d9Z
2AL/96ZU6kNQf0xVdrItgchL7/1sNBtmsQO6hc+i3s8gR7jcL2pmh4dv8r19N3SbDrKlhtRoOOso
CTvBHnG4eRC478tq6KbH/NwVtEH1yLTKVcV+klL2I0Qfjspuqfu38+puJqemgC/aCbKQO4sUK8zV
EPYOlPykTIBz2H3hhna6wThljVsq+tKe5ZYrQEbT1zydA7Pdfgj6x0ZgITRckZ8NWxPRun+t7/hu
0p1YosdSXZC4JubzF2nN3ySnVQfB8HEy8FzBbGOsMMhMmt1IcCg5PkF18JMvqalSYR6+azxJMRfz
9l/B9BkXsXJE9a0SzpQ+In4T+H5Bd+NCA3HyZzL0+xCrfd9GGomzmHKcRMwVDEB8oMPL/YEyWzfp
cF1uhk1pijaLdKER6es9KDEPnXiDJ89L8lAPdh2RJ9V3rlfkbfR/zVScAnsP7CgnegNGx41q05Qo
7oVDM2KfY4ciZzOOX7alWiOWnUu9j/XW9qbmr5CpGgrwccXkz9PaquishkCH/dslzl/mXBVDY0rq
yiKY5KRkLePTlSLomE4Yu0LGQlklo7O8+TmNLiLpyiuFxeZG5okowVJlSRnQSRBmKbzpP0k/jxqZ
pm+9UejMCJX9hQtEBW0s+hwSoqCRNYw7HdJcoBx8xJqytQk9BfsVwCQqYCxu7t3DSmv1fUTpYagk
zOVnladkviKnxozOxor1yfjJS9AE96uxWi71Wa8udIXx+kW0q7gCnOljhXJAAN02gJrsWAMdQPlv
K4N1uficmCqll16Vrbg+qRbp4pO2xDDLEO7TjkYKE1wQ5RmZbe/4/kO+hHkxk+A14w1bGcls0Jql
vdWUcKvQZu2kYI9n2ob3a/1kwwryPFjH3SRK2O6I3J3eg6jsRSxqSnF0ngmUgAVKUIC4OjbkXjQQ
O2euKb7TSDS4Whed5d6BrmmT84pTonyPWgTjC/3Ot47ur/CSKa4aSLC/t8QGmKQ42gb4mnRmJgsZ
MMmmBwDrnF17TEdglJAgvpMWmBo+/gAVO1lpHDvTyyWU6+DjCjHK5hrR7cWs9ys6D/4SJTXK3Ind
xeqvq8DM5k7dS+/g2GPJXoYYkrz1WhsoZD+AF15pHuws/Q0NBZmssksYNf9r0GlQdZ799uNEQVsM
Vgz+jBPccPB0Trd6ifX+XKIZDirt4CTkK1htoQCyKBnj8FrODHGpswT64p4znc6prz6D051Ypqzu
90kKVYif3mBkRmbsvxar1XZRkfNO3ByMv5Unk3L8c5P9PBnvwHrGZ/VxusQF8EjghOn9ECAVzVcp
MBgVYZPfFOJhaUSXytR8xreQt/e0EarGvDffHR3XbqVy2I3z+gCJQSSZnm2QULHIn3+S8kaP0J/9
VzXBIbA7fgCeH0qJUwlyLFtC0zeIPgfRPz4fpXXuJl28Pe8rzHy2JLoygHlzODCZpyHahW8FndFO
zW6Fa00mHApuppK5cWyZ6irhje9mx4iebMK67fx33cCSF5Uz5zQ93Qb0+BSHMVPGXxw8eqvuKm9S
yd6y0A+kmQrO7KY5UKy8x3ElF1UeZuz7aE6Q4TuT4Ot5ymRazXzDTF7a7FFIM+rfcc17VncUXg3A
uH8Mbe5f+L8edxov96Y5kJwCSTy8V6Fvn8uOb4wUo3s7ud9lMZGmfbLjEmK41+jGJcHDtgMzANI0
56NyYuJwhMCHs2Eu2UMKTQHFBU9xUFLo69JZeEFfjxo6TkqsWLHVN8ndXPHrZ9so7dPA59V+64dA
NRbnDmq15P1GBYleLx6uYf3zu8uYHSRLws4L1VKM+5q2qJy60ovXsttuQTrdyrTh7rZpwfrFMYR8
kHRVd0aA9mRJnBt5OA25PQAV4mc2q61WBRLs0CQC7UPH+uL+uakirfSR9WsUxfkZ01MwW39Xqel5
0z9M+QYPK+t3sfOYo8cIBtC5jDxmP05WSdg07fL0PI71kt34Xxz9j2EWhQNbKN0IQyo8LFTR0I/f
K9iNon7J+M4MFvNPyMn2vRLcSZLMt7YQacpTgJ9w0kp7KZ2c0Nm1ZwU8yIk1D9rXi0SPS3atJ1mH
aDoRzmN/s79iNIpQTEYlId7Pb6+EEcCyOrGtpC5GcdWOx2yeQpeqCr4FhtsZKOOoCl92gbp8Kc7t
lRlqn9t4XRqpX19xD4Xp84Pc/ZSlLM57YyXv2C6SFfVw19aC7P5uTTbculjs3UyBGfBc8sOR2HXD
f/zNvMUhqUL7sIVhTU2Nzi6SGbpjfCsB5lJEsj3vQy5DfTC1y/E9QZPhSwjz+a+U/Of1zbkn1TpY
q7qZa9w5I342lFFU8pBQ/8uZoHPALGySUhyTT7Dlr+4ely9miGlA9AD4ruIHEv8LBkMVNx/lFJw0
rXgPorxY4qTcSE6w5FCoSeNmqt/g8Af8brTM00zlpyScLli4f006IZ6jZkLz821TnvoWkxs39ECi
C8RmZxDXLKdphlzoLgIio93YeXWWwtv0hOSt3ydW8McvBx5+CW6bRulqJuLtEPGi56/TxM7GIysU
jtexxVVZkhVyj0DKq/9uxlAO4zcICcr3x3UlkLt7G2WheIvOZJABuKCWZRwITBu3WynAKl8LPwfu
5xifGCgupmVnvPNQPlzDDGok8rSvYCGoCV8mQvi21q0VwKeNdebyeI45Ev5rfvG8WPSZ4YRMAOqu
jJ5Zfp1ST8smyyh5nwH9Vu7aznM/Jkavmghc6u97oPVxQIOvQksp/buxoJQ2Hyyg/ygh0l7ML5tI
Ccs/S2wjWb422akPTnDh5NexgM+M7cvAtsx3N7VnxSu82POQEbI4dfrw5dyAvr9BOofgYK9gHvFS
7cl427VYXAZrTFxof1SJTJj0nHmlQo4JFQZas5Y1WoUUl/ppdClYARo4FAonAWktYDb1Bt4nolCK
5x/iKZM7lb1+H+3vJxrdnN+AkcKRF/27tppQbuNwfdXw80vd4Kp36yuhByl5aqsk0INrOjUyLNax
yTNKviicxpZ4jZw0vBQM2BLPcKjFb6BF515/IjF/LnYok0+NNU1qABnlFqEp5BDTgVSSD1L/ikNS
E7oDZ9gLtoDbFsafT5y7CpE4pcuboi19ZDCi31AtAjK1U+n/OBINwLq1f026YQbKVsEeH0BkoKcd
zfMEICd64s02yFo97UzDPsNbFpmUrELEcgrbtMUuNPPWQhLo7rccqSKsHybgqWql7bnWR88FEVig
bisi1e2n94WQRT1eho1WafsM6Hj250TgorJoD18s/4dEtK/LUfWBat4xxmq+nPtfZd2jILoeheIu
+Fk6jD6ZaqaoDWrt04H40Jc+7FhDFXC85V/U+znPNMKLjcyhDqcjYGprzJsyHO8s787BqJ6s/3IL
Uf8uALs8nz9daBr0xp5xECKG4MDUoNSxCk9+Byom5Oy8o/E3himO7W5XWXe2DaTDbEQhM4V4OOTZ
pNmwxfe4Pjh4QlCFKqddgy3QcMtjkKqcXSWlj9pjyCq9pu1V4tCfl3RoqcZb3ubhU1vRo8tZ4q5b
THQDQvFkU9Xrh72qQ0T0+eAKyd0yQMejYq7gjLd/MlvPJD02Lx659JvCoKXR6ENa2266mM5aa3of
A9sie5sKJEVEmI5vy9MAalnaWRiDGAn12luLCd06L4RkGpdbefbLR9Ennn1o37zhPrtS011fshvi
4NUAuASAdTvqjKrt2Lgmzb9h+ocwrdu6k/1K/ExoCHrt5GAX5ruigB1WaRMUNfYagQyj0+QhYfPk
dI3IDPXTRupnYsg80Ww9L4hkRM47gldDqMDbYNbxvfYZu3W5JwMJAhE/isRlYSULHwFpLGclC4bp
dpz6dSOf0HsGxEkjrAp6Xd9KPC2JHuHmANouR+QKt7kFHTxSOx182JRoZYDqKddRXX2gqxEqXdp0
YL1UNIQPcDEkJpQhNTJDcXVNptjG8PZN4UzAHjDdTpHcSaSTLosuRTyor85d4yVq6jh7aSk+yjIV
5mWpPx7ZqwIUdNWP1CCdE6eo5A3qzDsOKtJAjfR1C/vEuWZdi/px7uiZtxJ5R2IGoQvrgHtpJoTn
3PnfePLhQs4ZLTPiUIVscSkWIs0O7DieM+Obx03p4kd7EMak25ZxUnsHAa4IXbRmtdmXiTb/Qg4I
lTYeMQqqzVrHA92k/xOImzcRqCZrAELz7prwMFE9u7gAw/HMRmpdSLkMNcIj4YX1+e1bh8OGUx9N
Ypc/UzmohnAWxtimRFI4ppbJRJhCkEMZm/UeyYERphyssWKbfAjlJr2BCnIQlXa93tObUK+2a9ua
onv3RyRkg79CJqAiGw+nuZPDdKhttEp6arWtVrSK5yipCsQsuFps/MFYp1lxZ3kW0wqruc9bIfse
4wmz3dqz3eNHuVgHrwvmf0K3yIcHhqRr1A1OkYMOBm2uavmSwFRTbw9yugaS0t3CoozqMC61v5JF
BFZBKQ8hUKlUbKDO9a9tGA6Mkqll+aqyHQ0PKvlV1rL5M8WC9bFqMF3wy5nosnzRkVaHjnby8SIv
zjJnydSi9qQPy45cky5ZW9kQfnwPuMMqIJhXWnS4OfcyU4WeW05wwEg1Vib8Z6AZxj5PCDD1yi+M
9tNAf85iZ3NfnpLXTCie8gg1ywrWrFbpq/M8syTryDgsUFkHHTwlx8vQDA/StPaOGU2bNvKMMNga
0ewMLew7f6qRJJ8nLhqrB7X18ZMwW3kf+ebH5Fd3GHT0gbHp3DapBhRiPX9+S0rfBjwS6R7Ljdfs
zgXciZcBw1sDKvwPJq6B+4PEjUfSTVZ6xMbuwWbh3HzzkvcABnxNV3h8sdpkIgi9xIzCP0xCtVnT
oHTia9xjgsdAbiLOTd981/f1K/uMUM1XyMJ6x+PV37Lp11N3ahFvPKPBY8lBrEGIs1atAp7Fb0Iq
1cEvLDQmmJkbj7Y+dvvY3NJmuJ43HrbPklDKs9EiQ5s5Ny8UJAq+swDnPYgCve/NlYeGy8E7IN7c
H/Ak/hewiRw9RnOnuf+V7i+NLjlHHWcvVkTFrUTmAlpR/Maw26TuA+XfAS/YxFMjW6IYb37gI5UG
OFCI1mKqQBpj2+O+RptuE2GFxqtccyBgsHvElzXW/Ur4RC3ccXw/C8tEi7D5eM2umFUjU/7Nro7D
ZO0evj/JO8m4nYqcxz3YDy7d2KRD8PmASTUbGsd6rsgudy37mNbVljrNXMlgCzjtabNyLaIfaSGT
EeR1z0X9B+XdVXKDWQkQr7LTYMq29HO3ZO2C7wlu8EODBaXukvKxkbzaex5i9KKgs0xhG/1WH9TI
BP3miv34kjOmJ/hDy0C5xZmBwfdDfi8pgKwROKyJLfVtwQZDdha3CrFdH+3+PE+6Me9ikz8vriI7
PkxrNtUM1zBlWMASKOhXHWbeR7UnkA00TopHn/yo7xZopUBhDETUgtpBGBE9xhsIqTO6c1pL0hwR
WqwHOZsFSLR+oEpsk0HyFmuCIlIwyuXK/R0z9V1rQdD6x1RHMFEOG7327STCFV46J/m0w81NwO5H
KKmd/0fJqVbgW5O4rjDw8s+ijxbYkxOtRxoUuwFIRJB36kW9otyehGoG7lozoW5qnlrFl7EVSwwC
CXZdrEda0eYltcsZI11Q2r6/dGjRLEbu23cIclIlpEQPTijLt7P26B693VgWtFfb9Jd0bX5amHSc
QRpsJy32PboYuXxgAL8rr6SZAG4Q5jIXSoFj3MWjJSA343YsF/EeirarHxeKmrVuNeACcfPPMHBV
Sc0mmQ1TLPAf0kHe1RQU1m+JX9+HIS/8xgx8BhGTEPXDSMENHteSzBPw3KDjrGrp+HEQ13qOWZb8
r8rmmyNo2dAF3s4ud5y9ay7fp8rGEGCBxBOe4b765qciWve9G4vepvl7iqDma1Oyl7PxU8dTV2Ep
wP1zE4LcEaRs3GQZPAWWLdTtW0Q3ts9OG5DNeawLWuW2CcMscW7HTSw9evvJUCAj6qZn+ZXo/7tl
nkkRTy/cqJU66NR9pSKM+0uibIpxv27M//owTOZ4HAHKxtlXZ1veKm92hH9OQpyxK/nK91byY0XV
RPEF9frpVjLrzKPGD2LO8GAZqwLLAzGuI6sDO8FsOqEnRRRSg0+CCxW3E+V/Hl95uZBWJUCQea8I
g+RnvatynROEkn/NILZDTsJ8wYgJkkw+koGksEQzfeb9dCUVNpy9sVhopJzH79Af6kdzsMbHWpqV
SwZOjSiLUKHMldULHuce8W2icZ8nnkMwKkF2Nkvp9oA8B5/ggFJz3VizyTjW5WB1UX1QkOmeKGoR
mkWeyNnyvHKY7MmnfkASPcDp1WZWBTbVRARbt8rZV7av8x2ayHIlQlQuILc41KUJ++0orsDbtDCE
hNiY+fW8F160U5nxLtKAxBON2EZH0i1ijv/9pOx03fJDXMKXfS5rHlhAnI1cMdaWkwCtfa1B0Lc/
MMknFmGrJRnqkwJc2pvUHBvRdsc/mcVsh2izXtMfoTKwCpBHoY5Oo488TMaEgtYrM5xTidiL36Ks
WS36RZe0b2SXg1eT6p7F9aEezBxRrhxyzVMIJtNjwqQS1HDZlnoS/JYUEWLMt9MyluqYfFSl6TUH
/QzwfyHv6lZmjs8UObOZdHx8zTwhIATFqqqQwdAJAC/Z+jEqxK5X1JkBSkAL2xvL9BUOJlY3j5gj
SUZJCClpZIjoZOrmKuGK0Xn2xxGi6unXYoGYzU02jm5y0xJUetr7ZmbSCL0hpCgJz+cWrLDyksSJ
pKsRe0DGU+Whbr7/F/kA3wxi9+2bvI0VpOWHKqw4qGbW9a0wRrmG+XCVjDpeNTBw/zTLGL/EG8EP
TLn6wC3bq0AcqZlp9OQJ50N724c1RXEfjXG25QH9p2xJojpp5RgIuLU346scAr10MDT4uj/bLxqO
3aufZsV6Abo8EZz1rMXb7/dCL/DCg8zFPB//5G6sgNWXI5+qo6EvUBcBIzb+NJlvKqMFBFqJx0+l
NVpBDs7uxvE5QYwW44Tuz89Zop/CfNftcUd5+FpJ6UmSb93U8gJtZHoXifmwEJuEM9Kt01xVt5d3
Ut8PO2vD8gSHiR2GPlDXibAXwBPdQRPfzt3HUtPql6DrHxDB/+q0jekFnbTQK4DFM0YANlJ2PGon
VxIyMbu489Q9lK87uyaiyFB18gsOSun2wpkQxLhefMDbev59+ey/W5kzazcPq0WrDwiIHcwJqCE4
jqyohAum3WkYMTz7fsHP8xWMb6+Xc4smho+LdP4M/x2eK7d/17F7JucHxuQb3XOqRnuPj9+zPxf6
6bJEoEEvVPCaY0n++VaYw9Nu2uQ6omP77v7nsCCz+HwXEaW3IVglKFN8oKb73Fj0KS7snw78ikYO
mF1RIQz5xcUphhZphsDiMibZWf/QiyARPUvDJ6c6Faioa8JVTt+99pTsOHYGmCfwe71fIREx6kgY
FZ2HqyifKwjohjPCemdFTIKOD7rCDhUjhGnmKo/4ryzwX1J0r7kjqjLf7lhMZOe/5FdilQn6v5kA
TJIWNU5S0qie/zrHc1v/jeK8xFa8X0/Izure/9670FSRbBxd5sE46O2Hui4W8aivz33y0ga9O65i
86xwt+BplXryG0hK+GPtI3Wl6DGfINzI2Z5iZzdB1ww77NCWf9oT4ZMKU2bWgqvtug8TPvXpBE0G
VGTpMfhByPWgPpATIuPCffWzdhfy+KhMlZnNlNWTGMPcxaZ2v4nLBYml10j50hCT0ztjgzFEV96F
oRO5TKIfe4z4GBwqBPDm/OL+RbIXpACcne73OiS4gDK4TIunsdhbTpqZ0xH52X7brEZ2vbIVvie/
g7BD07B5JpAa3EbgkClOkUPCt8NGYClPW9VtlkWXylfou2huYs6jeQ+NsTDStMmQGLfQZgHkZiZH
S3diVfZxzXN6XOE5CPxP59Wak73quMV6EVXsZrkmKKxelT3TI6dXkZQW9yDtpNci5s71CvWE8g8z
mqE07xmLON3dZAGYioTxqQEyN8d/dOPkYKrPRjoRIdjRv1aWcMXJaz/NPTga6sl8LRDxtkNcIKs+
ItxllfwqoCU4gZuzbWSYcK0Qvg46+YwqgcVdjshLjUI1zjzQsqbGOa0ptgQ90zqp1rFehbA/qsWB
+YJLHI6iprNXR7xIp0Q71LeekOHfjmsHsk97bxBvI55iatIpFEztcFy1R3YtyFDyMxn4e4hxmihJ
0H+EwgSh+WZtzmosLJCpdAXNeAsdKMyIZSIoVgeLuRWulOQpaYT2A6hrGUVE5f/PNpBnDhquB1us
RFl1CcrdlEWDi0mdqXxmoUlm89CTecmtkHrPMsr5f1g+XlrIf33Jg7BzQ70/H8gH783z8BAzZlnJ
coPct5m8K+MDRokDSx5/WubrzmrBtDm5gnNm08/CUZb8E5GowMBxCi2FY64xh+Jk0LrU/xPgJyKg
TXLx5NxJeL/3vrDRK2x4AQOEGqcuREWm86Q3DwRysqoJscnlUhoZSzmC3ddUlTP5PfcatbGIxag7
6sCklN3/0ZuHEyBCpdDXqGcXz5wQHb91M4OfRFwXvwTmqwrf1Gf6KN9+mS8CS/kJRhSNitoMZh9R
LwiylbopFvQMn8MUL2PfHIyETcuYVZH2Kd6lwt9GmdTrvoV4EK0NleJS0NF8la3WZnhj+8v2UcP1
XnmwWSQ1cjCXKQLXcoeuO1wBfILT55ZlSoQxRbHrK2JnezbM8NPnVOm0ESY2jx0MCShe3qUE9b4V
wL5W+NqQZuxbHoeUz/obicVwtMiI2xDlRiMO7G/zjRBeGSGXCWtRkxA6ME2ujKFBTZlBAimvOSlX
WxObIFMrnl1xRI8gSJ75o6TqaFmGEIohZazbQhOXevs1nWTRusLGaKcTjB9L6a8L2dUF+qNPb1fM
CsSWS3U0agGqN/g4ek3PJXrZpoE03bB4u0uMweeGcvNQCgkKak2FqJXYTtxbFz0/aQZC+EVRWJFx
FiFPqA7RfoXnZArZOIz8r7zVJ5vMSzVgqVxCpYFirU7fWCWysJrhARqcHTjBsTmw+Pr51+uzMZQf
Q4Ey6G9/hCnq8+hAHr4w0q3LdBfdSOFTXAeYsES+w/nGD7guwi28urB5f/CeX0hbWtn7EKsKAviV
Q2piQwAcKEgi//bk7kCGbuzCCHcaSv7xSJXxGKEbmBdB+8g6d3kplpQk8n7n9m0WqNLkHxcjgyUB
EqOp51TZgP0UwhdEDai52xKwTDFOzRgxcSAieGoclWn7J0tciW4iacrW2gK1JUe4Grn9mTrUbDrK
UpQopwQOa88qS6HRGzqTN5jtvbD8b1TCdrSqY0ISUQZLZIOdJ05qgg+ZbFmsPxc93Mx98vJ5gVzr
umdyXj4OkA72EhBauKEvqtCu8JRpz6pmt3Mxp+bSQLGjvfbX4bA6ZoeOgnp0iOJLDltbOH4pmqn3
s5sLFSv+3sqw3XPWgbDSD1LavvOhuOg5OvT5dojRfWUXeKkojdgnF/WH8ImrGiiuSW8hsHuX2QSQ
MiHhbtNEcf5NBGH9MOjQDtY2cCnf91jEVGJTuPtLgJSF5i+9leTvh6t4RMzau/xmiGb9jr5udGxr
dd3XscuciqWWBdrgOQfdI98fCpiUVbXgiWdIxyI78KWUoeT7AI3Ak7HMKQ7A9hV2YRwJAaAo6Ej4
WAU1nmtOZrYzQXk0iRUOLUjn7KQ1NLIPaU3hlj8oYcpahhdTMqW6nEPqJa3mymHWWP7bWiBpdCYA
iwIkkEb3JjPxP+phVc3IGHBic7qF7ESBEBxu/Qwrul7DOwBzZPtuqBRS5AKIgV188gRkJDYQrmmB
a9Q7QgLG3APfhTSkMwKp0S7v1FndQYEFnNAWgrd7vQzk/Wowlk0a77+y7iMrBZNhgfWi3us9KaL/
m7hQrZtpvTxufE4um6ZspsIOFpwbcflMJ8r2KHP5wXlYqx27UBmBKVyWCOsXPC7FBMjULnZfBQZW
UwZ0xEKz9G25H4oDcFU/5uPJAfxe/6156Gvhgx1oCLx0H9/bMaft+tyzb8ghiZEkOxGg/+/C/rUP
lqpktZYV0ARRjM7cfodDX/48wiqnBCMP8BhHkH1E79q6MWskK9FDf8U5t6GDm5zQ2k8uMdlyC/ac
1wB03L0sIReWDvATZUoJAHJebLKqbWGb22ZtjFkaC+X3pXzl81lT7UdWyt7ykRS4jEZvVGvKFvzw
NiQELz2FbYSD3V3dalLA/skD8rtxoNC2EBXFOxH10Nnknm+2jd/QldZh6VGO/4/VXJ+z5auMZoh+
YBA7xSpNN7/3qZR7mCAV/tGlly8TRTa8yKZB1PLZj7Vv1QZpmN5F4KKcfdIMbpIDOcb01vL/QNvm
2uX3OOp6iNSwu1t1ZtmX5l9cuzK9Ce4zfMoSoURFbrCowSxRlvUdGe6LgJ2/mbx9KqEszhpklxkd
zJSJB+CBjV+ZgiOtI2y8dsPTqxoXVKUzMkSYm4N+ru6F/AYd+AQh4YLOQFsRydCenbzXqxHJr2aD
1xFIn1EinioohpFcJzOCAWGuUDJbBvU1LApLXNlm5GVg6aHNg4Hd+n1TyQY3e9bv5JcCkpbOs5x5
XoEmr+omkXxovXiz93PuW3ZxkBhkBF8AucS6nnz60Hp1HgR3jjlC4Qzy7zvZ2sUiGAfA8hjPUluS
7ydb0/8UzhEcdT7w5LpYgNriKZnRzGbJGBT6vYWRS3vUGan9x2D3BYseMSBQNdOvO0+WpbCH6n8b
6MvtQvhYZR94n0k+L4XO6xVgWjCXZqyn0seU2iQePw0M9aqOA9cGzx/T6QEF1F4esYOWeY9R9MdI
qsArE/DvqN4/wL7HqAMb7QqcXK0UuEjjLX6f4pdikaoGaiJJS0jwOOnR/2i4ALI2VIhZZ30CYOFO
aTyvEJERKkk/fh4sndAM++ONhNlLMAOY03iGgg4eea3i3CE7ts1+h9BVGoai+TuaBjR/eMmgNaLB
qUO6hhHUn7T9WP2OxyyvHloUzfGCzYK+VYSX66YgzJznOP/55g9mrbMap7kbCOA8JepQlS6jnFcb
zcS8ESCG/lk70HiG6Y3gz/U+RdtXgh5U5hTACs9N3Fs6eSlgMdYm/XMWBANUN3eApFLAjkJPdsWL
gZXkzefWhQXPKb85xSoPNf1Bzhw0IqM3H3mQNd+wwQLikNf6I7o/3enu36/R5G2fCrr+9fVM/HEo
OBhigHfVzHaIqXZ+krY084xYvht5z4DaBO8L/5pCwZR5mYmxBJjNj6meG6p5q76V+qRSCddqioaC
dsY9yFqXW5QodaTZzqbfQ/Meqt/oT9CBfFyQzB7eLrMPjmJxZQfNyoPhYMGTy1/qWlzcU+pqdIFQ
5/a8QoEUBej267PZf+5Ixa8Ada3EnTAtDWIIFKojNg709ZrGX8bnTQ/XfN7zO0RQEJB3LCNNYLsQ
Hrqq5eTvri2JdsJaVb+tgmu2q5SEIxyvM6o8eWYgfLtP3oQYiwCYD9bYw1REQyAYKQIvbtcc3Pyg
zgzHqhPEfXQ8MDlMzgvHXoSCyy6RMc7TVslDM+qYaXMWiMLfhvKjIcHY4j9zyFxZrzz0aZ+GmZ+j
YiKgcuZsUUOpDFz/a/ZwoN131xBapvQdhnrF6Nd7jA0S3aOIlySAO1woDeAit/IUPTe+UZFCPVce
upm0gyk+Y6mmM8HYpdYfarvwn++pccum1uMUmT8PMutLeFtRkZ0rRt/qxMbDZ6gzozOkn9/gwnCp
H5230HS23BSXOSYxs5HOZgixcR55MplG6RZKGEAk3pEGhumOqdHd8KvC8F7mpxZfmxJwrIFRkV49
DVILtZxTUpKtL7owK/t1GafCvbjRdXuZTaJkbY97r/Ag5WdRV/tz76eBT2g4yvzEUlkXJ5aCv2+/
OGMRYMU+IaCA8s2v03CMipc1N5OnfNi8+zhyC4wv8fmo8E7f8/zJUifeeM5hVM5K/YGWCHapAtdX
9qoH49XYP7A5cirsZGEOl6GPFBoi1tswy4toS0+nckz8n3sbBqfD/UioWdTMs2NGX1sNJtp8huam
fWJJXHkoXzpirg8oD8GMB8Z+pFqr+ZM704j9dBtStRgoLO/hlMBRm0EXwVgg459bDG1uH+zXlHgM
fJ19Ux5KKU/M9Tw/MCRQp8g87uug/DEKda98G1Sb+A+KPM1BScYEdHsypWrss+xt7u5ej5VArMEt
pyfT18d4qF7r9VXUn3hfl0S2Cxo//LFUXnKhdr/M3VlIW6avH2bXgu0ppKgUZ8Sa4Q0APMCaEVyf
gjnjk1krPraX6md4P3ebkCqXPuMXuN/SlrqAYyxv8V8iJRaJVxJJSpNQ9oblG4co7inaDyIxm1Pj
EGnX0drLTE1Dw5hSoLEVxvbBj6iiI5/8bXzpddjZ1JXHYs9IE7h17ilj0sJ4t5DnpexM65DXOcCS
jvbMXQloU625hRPV0vY4QNVxK1oxjx3a7TcWxriF4zXWkLkIAFkXoZJzryR7ZfSTvRHzss+E4efw
b3WZfcsRR+Sf1UeJ94HU+h4YyNQRl358/ol0R+ekjqOY2LbUTrPxlTR16Hhyv0KG6AxExNe6dRS0
dabba3BSubhg5riQhokbApZeTbhI8wb00Z5x5hCQogEHRMcSTpDARixaqPGzkB4zFJUGGPRYq0uS
43lRVH0EmhOmsIq89jpbxo8SPXCNDD0JNn5db21s0Q6YCmmmg43d0ZqES0U32GC2WkF3fHNnYRkD
Dw48eM4+n0Es7f72VCNTMDtcHZPvNN2b4Bb+1SjruLm/WHykZocFjh/vqpH+AJJQT151Fjq6YXgi
ta34zH/vwHZm2I7kqtV8NZ5Ztus21/HHNyI0Z19KI1F1M0ggOEkEjlcOM9UQijtC+JM4shwEuwg1
c9q69n3nXegDjP6rIetoVPpbkJvG8QbeVpr7HnBIq/F6tOI1pv8gVZJfKXCnAr2EJ1J81ATFdHIY
KHqWebrkyn0iLvPn2eU0KvWl5DT9vUmMTCQI+9rNmhoK1Yq4z5ywClo2taD2DuvO5iFkpBAd9t/Z
qaECrIecyA+ugdQ13PQteIWkgp+7uRRhHo+ulf+a/kOZL0VtCjnbODhbPLV2+uKSQhDaED8HH2f7
zvpBFBUMW3If1Wdxzwb9Mkfy3718p/xoqX3AFwKwsePr3LHAWhZVgWiBv7bhW2GCFGjYVmf2XkpT
TWG/+XRl0Kx2dHXItKvrGszRhMVqqvgMy0p4Mea2iqoLyLHyKPPU/6pCRS0c6fokc5AWPyCWUCNn
SPRylWjGkN0GX9HVh0g+rYTyEoB8rlv8AIizMzjk3kACQ0mw15xWK3EPj3ln4x6ZrMvWhNaHbHEf
hLG8tF/0ttyMOJ2CNEwLYhkYmdRXUIYzT2uZ6KLOUGoS5OCgPVAXdtlQnQlkoFPHm6EM0oxayucn
DUkUNGw2zs08KUoRJUJjLGO5ie2/1FDOKMjv74w+NyM0zh4H5BqWGjAKOIlF0ZHxiy+PjJBngIEx
sAMciBnGglYSTkK77PmqMOb8yIXpkm332v9QjAgGvW4XqPMmntq1+nChmsqdg4MHw6mtOVJTT/hS
ISfeLa6qZclFcMv/i1g7iRLHXJgruXMf6FX/0NYeM81JVymoYU3uShjgQVzXl6N6nHx0jgemRzvX
gpluU5ul+YLdBeoPyThGxbWc1qeSLkp+Dw5JKNTutVPNmhixnsVT0gW2w8849mymChGKOUYrwipM
y3NqBCJFXn0iaM7Mhu/8bo3wfJpiLVbdDpJVwWXqq4hDXFVoiJAkgsiRhyI8fet2vDo5yT7gduFU
Dcn1cpxbBxjIDzc1QTTmb0jFVAPrb0jQIIinO+HvzYS1M0tI65qIm+NM6GTefCtp9XiomOS+EXUg
io+R3qrD7BiwHJIn3mmZKOOTrw8P3kqFbORz8q7kEHdNcxzcLKUjrHrpludkabKsC0DjNYJTImkL
YzXRpBDwYK+oqiyYviL+9/14kZT9xsi4lvPeToGKQVq7EjGpC3loIc4GNiKv2vR+O2yTqXOmXSXy
8hIi/HgsocaSpY2+ZpaqVXRWbxBj8hbg7gP0e4lO4LmcFJccXIJwJDsEO/swGpqK2OSmYeGTGvTR
GPFLODteW+inFC5e2msDclP+R3pwuSb24qW+St/hKmqeuEnwjXEb8wkGC9DBYFtEApvB7xZ46Tj2
LZSiusOzNX/a4/2JqXviZRtBinNRbqSHJFTg8oakrDCN6ktW4UDjJv72tT/wgJh5U1FA1wrF8/IJ
d/nQcIb2c41z6dRUOIwZAIG3SvP5fVvAUa5Dsxuk4apFzTlJAoC4HqBJe8SMbxangXGbQQY6nsdz
C/aQbzw9WWxDj1+uywNUwBEYMvEWC9QAQ5gWZlGLgkCjPLprHqv292tvOUov8Y8Smxtk+yJWB6/a
6FoDPYaAdsFDxDDUeqoH02yAf7CEkGq010U58DfyrowQqNoomZptSpZbc04tOiAnhUL8t/8HBBpl
w5x45KXRXCyOV8cptyCJN5Wf9XNpNJ6uwshTzg4GvRArcuUL2VHaJ79pY2x/lVtTLXEHRCrw96aE
Q/Uv4rTxMP+en+Omiu/cUJ7L2FHhB3m2odGP7UupPMXyKWUtFHlTfRCXjjj+CAI3x9nUqkaM0+8s
dmamOcYGnxBndXFja/WNe91Dbx7sIK8dRhEpwfpV/PwF+5+tG6VFXzprCzmxYe1DsAM5dhjJMiB3
wKvVZMbeV85Qj8jmPgFA1FGX58LX9rJLjY7tY8fp28Of0Jvt2hGVcrgjTPelkQsaxI4sE14J8Ky1
vzfzENdoW0A99tbo2RCVU6SFP15riXDqiEIuxHdtPoPTr7hdVxyGWRuLsqpqdoNTE31kVYNXk//k
TrdESSkedzizFUk3bKF3qeRSmx10UpJ5pm4FKaiAJpGpw8jgxWdesZhYC4wtDvu0RDuC7Agv5nTT
fskT5Rt9hErmklcwXt/211SztJDG8wfws7xmdVvD00RiqyKrRXr3yPLoIRUCsp9qrQD2jikv+w2W
BT7MZ0udjjqwW+mVfpeVRlwP+t2xmURk3TxYouNKSFpntxHzTT5eRLWn+TL8hTaUfUeh7aCo6yBp
PoBVJVDiwmFzZfH9qaGxSfKASIQ+TRNGxrlaj7vfuZ5mMSKbcEXCRhaP54sVTMdRgEJuyKjNiyh9
nKbEuHhvzhSeGSq0Hx43593B+0YEFh8PR5Voq4fT2urBIkcjcRxfBCGgN+4xCrZTMuyiuHlqPiss
/hok6BoChQkQEbtAkFIGVuYRdSUSKy074bWhxOx4hW6QI3sCH6RJuM4C5ElB0Djk3pvPpGi/nY2N
jewb5J1G/tY/s/Uk9jgJbMp+cmqJXlTHcU4barcGlDNumdDjQmJBkc9SW1GJ8nM5yjfGSbPGAlVh
ISjFdWN8mGUz0c1/Rj85qfYVlOsVRRZQJlt2ukDoOJf9TONnUcQgCjx6cR4jSOzqDTj5c7qdahnw
FujFBtXEcuw/hLQes9Zx6JwRUi/vgDhCTp1jMxshQBSBbNzO5EgRkma0XldVN9pP0mMl0G+ar5vJ
Piwkz6xnCSTM5lmPsqPGzAqCVlh7LNayke3VzA9F8FzHUAiycOBPaij7VLOEUYWq3YPzM2baKnsD
cLguVFsiJ25vt3QjP9ZwBx32IAkipng/6tQG5bahaRuoXiZZeDd2DZqnOD5nwHMczm+ZCFVx4gSs
8XT2DRzLdCHpCRb7jB9l0i8sM92QuZrj8z+2BlFviW/tHhbixivSzfiRhbDvKO79veBZlqLeIrDQ
1WisJ7k2XOOS+zRdegZ3VXs93MBCn8MhMP8NpLnbef1vf4K5NSCoVNE9GmA80EGnWO3q4oqMQ5Ze
ULHi0b3yNfXDDUItR/+eYgZQTB8q0+sYtSNcN4/hefPWm8n7EHvYF0MuQ1/f3t+A/Ob6bTeje7Xh
6ygJ85dNRSojY6tUDehkaygQ54p4jOZ+xfFWHFksjUkT3TDbIpw4haRyRK4KfQtqCBqwk4rwmVWC
Bracnghm+NpTfHlWh5CjFysViVj3UThv0iaO/pTGFVcZFakjPpR88dCRgo7XluOgTOKhC7ttPfWO
b8RJXEfnTB3pNorfPOClagDI2kJ4ipyfdr9qmVFL9N130g3guj/cCjzDdrjIXOaoU/qDnJ69nBic
V7bA3Y3V9XQLQTUB9lsNK63As/JB9rdUrFGKNqY2vdBhc2mxOr2aeeSoz4eQX9ssRZrQhYq+JarA
8xwF7URkfPWNZ+IQBH2RaUpA32PTbwKsD1F0vBbitlbLymxp+YOm0dvLZTVZGzBSvkPce5umVX/9
eIYKjWU9+yIyyrhlzgcyECq43/7vrtRXIZE9pxIU95RfUPeoqpTPjOkHJ56mmKq1WwtWIe8Cz4HG
Cg2yPtBxsYB1ICz+h0EjSJ6Q/jmaBTUFUxBnm8G4F6g0MbF/0wfvc811/RkoCJPJplcqklZom/PM
0q0AJBuTirusp8eK/eTxwX9NrKR3f/t/Tr34J6EuA8/8tqgxdwUp/wGWj1F2QcOdIB00PIGPh4HT
plyvZ2LOrD5XtBC6v057F/Ca+304Gm/X4vX+t4R1EePuQ4Yr2ABatplGZccKg0Hp8JHcoZ4LMBJv
kjd+D1CxygJ7vOUlLPj7u4YfBcsQGi8+bMZ+nVL6M5nvDEE8jwJRPAFwVK+c4Z19U8SZai02GsSQ
TGvNA3Vy2ZrEw7alqFAHZhhiWyvDLpFhVOfilVmvROMaM+usfFySuQBWI3oLYAVNtyUX6ksPRrnt
5efJ0WkoRxSLMaGnRRGJHoxEAawbN/fC022L0aixart4VU9B0vS6J2QutAQ8kvqOqL+cn94kv+Sn
Iq5XPlxTD3uj2Bqx/njl8NVWuNe/Rkrtn7L0drnsu3bZ3VEHiytjZXROuNwQaykBWUvtcil/lQW3
QD7Nu5zJgwjQn86H9lnRCjcp+AXeI/Ays6PxC4XoOqQONGraPdMsKJyYcC5BfptvETIyXavMeOG8
GRFULmDqSVvbZUpP12DiMwumgSET//7KB9ncNDRG98lxCGZuRRPlLO0dmccredGyjKK9O7XEm6AG
mz6mAoFE/QbOl3ccRTuiFF+i/LJ4zZlLRrNFHP1nQNuvDARPtZPi0oMDznHcCzdaWDYXVKpWMUNb
2UFO3SB1yeas/jiw0kTv1fZU+YgTvLuu95FLechG2fpQ9cgNeTbFQFtGd6LweOSqiayV0uAk/iZR
maPVXERDxaYsYbXFwF1ABfuOInJdkEcnu5P0jrjFop2pc2kwEh0mtPrayp+FZdx68w2B5+xPN468
33m1oCe5A3wqEie69/jPzC+vRgUMLxa5KVt461oxnyRGIQT9IyEwSM71PgMAL1/HJZiwCCUdJbGN
cN2JwImi89EPyqRiTORqwyLvB7G1JDw8Ac1D5AVOpb+EElcHS2V8o9smcegEdIIYEsQt7jfgUhUH
4/ba3EwlbNXsPTkBhIBr9fPVmB0tjkpjZsVHV4jFHMGOO2P8OANGSpyvNlI2cVYA00+FukZ1OevO
TZMyOxv05T6UBb3mDq4W1DfTx5IOTIDBB8FmJrOENHza8xoby7MxEN4TJFRyxjLdVcXNsAAZyuO8
IDA5JlaOZcr17gVMW0bpU4NeiR5aAMjyZ+gRCycxwxfzaZCVGXwherTOD9TJi5lsF6w+vTAE1+2a
REM6qVJKO5nwI/MpGZ6dMvfoRWLuQ36LrQ/mq6hL3xgEE4tC76REs6YIZUmFylIPyGxevP2ZSI2G
v5Qy/DLc1uN/glSQOLJRtnwMvoNoFSYVI+e009MsRR3dS86cw6/qy3hhIGTRRw/qy8CzgyMWg0rS
+JzjlF/8FWOtzHVXO4o379Ji908YCtR9g++1p7PUxXX/0uuhaXg9UnDS73gn1OzIKz9cqqGwTZB3
5BA7wvL5xeQsPOZagKlxs5CM51XyC2BIkrPcXJeXXI2nbmFdMGdPYuoDCfqBejsgLZSHTUSOeEeW
YBpGnJi8jpkeaaP2xu8T0fliz5md5+jh6tksN4KAN9dh6S+7bJ9l6O1VRpQw3aEe4/dUENCE6O+H
oIuNz7u0LrwYc6nVoOPU+rbitSOGyH1+pT213GSzw3hG79YFy0pwMGMzPCE8wXxif8cRmwIzU1jz
F7Wg4DuhU6oPJ5JsgEcfhqfbP2/RI5puctapOaqR2sfsavUwoHgseTnmXGCG2ls8xVXuAUA8fLKp
s6t//aVPt/ErNYuTpmqcgINp1afrhAiznTb5r+Tg27q151tGnA2gWCqPYTQEA6lk75yVMdR3YKmG
h0lFWldtzscwPklQE6SHk6T0zLj+PfA0Jo63lXmpRgtGalHTg1JmHvTqn8n/nFSWaQzj0ORGfBHx
GEVZ3IV88bRN6IWHvSedcX5htbRfHLzjNq/HG0dtj4ReOU3Hv4QT8MLWHa4LRsoYkELOuS/v8Nbm
c433WA1ek0+RkhxxHD9BIjaoPn448IZOz5FnK4ov/iASGc6BoMnDCbgbiBbXp3p9QEQccRG7HiwU
cuDc5JSkMD3S9ri2LpUfL2leISVRxu2xpC9Krsa+hhZO0V23+6uDo4vZQ1GQVtgf0GU446B1CruN
PwUrcfAkSrM7naJZGcn3FsYsVqVr12c9A0EXOytG4WXYxwBJj6mZ7Y/6jidpnN9PQBR5I7k0RO0T
R1AUZxJ8DCMEtVDXX3UiXMTpTY7y1Gxx2p2/jKzPZ55OSt/2+H3jbbz7VBuHma4u3PzznPXwL+k4
SqG8TLYvVzgrxE6PbGniYD0VkVMYt7woQavNU4EmJGItPN2cw2x0+pPk3+Q2NKS67ox2SOTNjBGe
2lqrrmQZQwyiVi2DsB3vsMnvZlHeg3k6vOnfQIvmZ54F2DqgQEbPhuxbjFZaf12SPV8VbxgwmTwR
T4ll0i1Ha78rp/5OB3OiCOWLWOPbOjiToEiuRk9WMa2BVlhOqhGeG1LvEEDPC8G5q6jF7gVd25ZG
K+LQ4G4dlknKKmXB5nlQb+OcfitRdXBTD0WH+HVfJ2bxwRjdbf5jMJd72k+heGrqs+S/mE6mZP/8
jqQmDAoqwtaAPh1eQs6PCrx3mCMVsuhw7RfQok2yZRAHqum5H6t1Jft9c8OW07csoBCb0x0wNe1p
8HlA47AXK1h9T6BRLzPUwls/Tg7l09zS9VvPRasq4mWVJ19+zT5zImTgzC0F6FVOwfJ0HSrxknK7
ExB9pluqfMs9B05TLs9RvakUy8LGzW8+hDDGHN2LgwQwYWPMQtoKv+akexV9x5DgmU+orWi2/QBV
0EyoH3VISm1jgWo8jwgJ+h9ZmN9/XHvqJDjcf4+9ZxZkWIoIRmLgbBBbXGSyVWjMl6xmrJlpfICK
uG/V0lmpQP5F5ZzBVrz3Sz+LNBQl+husSOOoueR6e1+UfmJ98ucjsTJiBwYC+S3dLlwFJESyFqbA
bMEvv/XQx9JdABhWTkqvn3l3r5krxkYRxEgby5aPpeQ3lVGX1Z12MUM2acHJ8XtXnqp80dWBwOdi
ca42yAEUPlUBreXAi0JQogeJYdu5FjvZqmwOnF83tdbxYB4HxFbv5fZNzuyiF5YIDf8OHFpKjmcX
kk4PJi4KocHgMuSc96gfCxXfyCoCpqizG7gjNYegzbba8ydY9JZOHekKI3UWBDmO4BAYC1qYGJtu
X3oyY3HaQY5hjfBgdiT2syb8N1+UV/8GHPakDCGQpumVZLVyqi+idNuoiPuJC+LweCukPQHNJ82m
lqj6RGud1STn53pAsnSe495ZDH/ghddt65z9OQpQ1wXbp4mSDqRXd0qHqHTQwrCIxOfcNAK8V3Jn
8ZVXpbWppYcKSDhO2dDh5wEwSCkpDtrpVwv5Lpw5pMl/vj0m1tk1xa1CElI7UCnhQn2uNzydpnQj
unRbj1GEclGZrcRERqA3IafkpfdWHuXKuMD4btTj46Fh1Fk6jic+UhqIoxUR7OnVvs1OZqQGbina
YReoxOK8v6H2uiZTR08Fc0WZGbQoKMnyc+Zmwgu+9BIEzyaCHEdJC2aYj0+wtt2BdhR2kbAQaZ9i
Q28bg/FI8lqFqOXBEZsMlLSA2W7qSrJoNq+ErB08Vn4aiAVub90GQiM35bFVTqf61X6dJBOkBw2P
FD38nozMMFRscFWoYoobsOPEjYxsqLJHStjRgjrkkn0hbcW+cpJk4BosRLxQvo0xxqAIZe46cYTs
W9RpIpva6PjxH6CxFfm1JK5mk2iFGRzrPf0e/kIFi75GQ9AYGJMvLgQY2e1irhDpNBjAGduYMl79
MLCL7YU+wrPWdlj3ci69dv4Qfvo9CTDeWO60V8IC2oCCxSHu2lbbRWzhJwRt2weIcgLaenzJRsQ+
8tTe1PSkzhQzzYwHNixDg3wfaodX7RGicvmrOoy6pU/mOX9HM3vl8oZFSOoVEY3A6U/YBc8kd3xm
IobvQSUU3DKxsxmuVyUevaQGulKdS3Q2KL5Op8zweSkZrJsqWBiPJ1pMrDMXx7muXEk/mZpfatg0
oZzA0ZbnS2EjSc+JTQT358Qte0DzgDOpgmlrJk89myzPte/fHXqdf8cV7q/N72RUu/eUEgbOOfOF
WcnmZnBbHjwjgmda4OVoXgVkyVFUxihIRJd+GhGzNE1kP7TU8BJUFnHydKBflGr2jZn9SLh0wmDL
7zaujc6SHbuvKngrp91UXK85K/U05UmRv8Jr7Cw9iqbiO1TvDdGW8RuJIye5KS5DU3jMtt192SL4
aAHWy1g26WLlfDUMuIfN71g4IWW9mUCtJRJakGAD5GcazwshfcK9c63SeWm7rrHmDoYh1Deqo9uE
tIxUfuGBEBluw22Nff6oLVNvRhDI1rmrWOWEjA7b/o8Udke7Qr4qVp4WKQsk3XrFvQHDfnNQ9hVX
VFZWmjD56HB/V+cYw4HEvyDHyq5wrfPUzZ0q64mqqHQ/CORLLVSAGOFaM29dcc95DWNBDm9PDjzU
Dypysa1LaM8YgzI/Ijcn1SATxdG5pAJwVjxydqWZ7YfEcl3yhQ+CB8LqMPNLrX5fBBlto0fiVdOU
bdtHyU5OuR+cA5Jr49s0oDd7RTMxHGSE/1gjwVxTjW9cCdO4V/WBaUrUEkuzi2bNp6mzKjorxmSt
BhOEhjn/gm6kZFG4D7n7vX+s+JiC4tpd9SpkGGulCubGOsaYBLtsBKrJOl/gyRfBbNuVK+TWXL4y
35zYd12duG4Kmx9PL2Z3redgXZKWOSf4PxFOWoPPTQ0fr5alywW3Y1L9yQ+fRe8mZTSQqg0sLFJP
3Qg3UkfqUg0CaKFv59a7s8SWQpx2k30HbJRPscCT8eVkk/kxSYag4Y8mjT+wO2x4HlTA3dPiLA8K
bpcHOg8kDySyMF8v1ZMNnexFS29RSYC3s79HhneV6i2HLhjRi0uxPwtanK182b2evXcCNtHglfv2
rbiOTK9zkaSCzG+yNgU3Ieer6HK/0nTk516NI47orx2vMBmbsX5myVls1TPdVy/NISK6HmSEcRBt
8xVcDUlgSDwS0aWQaGLPS+HoLzWeNkRu1yILImyNPWDLy6v2uFL5P/3r0zOH4T8fICSDH0COjQdi
vslyDVxhGrssmp+UPX8De2cIVZGQP5LpT14x5HF1nvGNSdZdq3Mb5zH9FkwIU1y/tK8t2ptdL/8c
p4I37SxAJWWGvRKFk+FK0AbuGcfXEYdeGZSJi1WVpvqwkrC+kkRxKTj44M8l0jcuvaGfG3qjzcpP
GZRr+j5nRZaVvT4GoNp7w9FovKNUciBDuQewaEOidTo8pfy9FniD53U4TaE1yvyO9O7PzL1145yW
elo/byRYWwBVV4PFTThYCnYhBh77PRu7GXpJQ7DHgX9rd3xOrD4r4cijPSf4XG9jYAfL0X682hQ+
skGurpIOwB7QjZmjdJnIG60kKx8G1/qgni9QWTAKN1kBXjilkOGc8tbOptFoKeu6w3nLKcs3LQRb
K9j7xJchhw7Sm8K47uJGccNGfTtjuKceJJMeoKdUIhB+/8oz1u0cR37GUoaq8J4bqZNJSRsHNGgg
QJ7vgunb0qPPf1vP0yNVjOp9XqbjclG6YoBwaB8IMdy7nHytAyr6nm9vf1kURaX2a47pfQzngC4S
vgR0AqVqumMWFOTqZanVDJDWz/dEgJp0KZbdPQTeQ+w0oXNW92kZiJRoMUrMTF/ix/T/sRC/qJ2f
5eLMuZ2oTVMKxbhhBqzsdva2hcL+awumliXwF5nXD5vFyyHbA5zVRar/x5ESgjzgoraCCLh/LCUZ
sZ0OwWSeFmzRovcOMV8aTh1RZ/vFnijcAEMDw7uhlGaMhN0DwBa8s/Zq3qEq7iUWCIzdM/KyDGZf
/sqxtJT6hQxnzF8DH0mLnALR9eTB6BYzgT4tcgB8bJoJWKwHlmaJQMOQ59gdZ3Wom7jhI1oSGlKL
/JweMr8P0/KKPwZsfMXw+k+T5gBbyYGGvVm6Lv7qmDUECThHtKiWu+199n6e5OL1GM+ZR9xsUfEN
Hc3vyYRzaOxCPaIH5iZbUb8fywZYlQitC0rYUvnd0ehKkiZsuVhA9f9m/qiYrFLImmVKFJHWP+Yl
qTLKPnKo5w9u/KKxsRMhsIbIVqXorJeMhvHLI3IrY+Uz4GbMO1z0vsGVqZaNmga4CJFC5tpqL9j9
U/UGgdGl3gmIDt33jW0f0l89fsAvlCQhUl/C4aR+nBSwlF1t587zWVBljm24Binil/aSiwAtvvlH
FRWtzQolZa3PHnGKF43FQ4C8+fac2kwoTx04nXxlUrawZMHShYAU0f+nWbhlIwuJGkSnmfVMM1RB
Bwbk/AzfWaqxml+rShIszOURNxHZl7KZjLZzM/GCGpgJdp+k2sY2bYvpugetgOZIPw2U0Id4nbqQ
IbLG5O6CC4Aen6Pk1K4jJP8OsQYqffsYFBp2x8u1WjqTMNuuswKAxtheTT4fD/S9D0eR1y3BgNWJ
AIHF8F5nc9mg9RAyX6/s3+7NO5pl4URWfNFqvSKZO7ivYy7j215YYXY465yPlfQe9zqEKuyP0PR1
lwxfoX98VFyi0wPn6Grlf9KdtzlRfudizB2lp4B3w2EnkrEWJccSw5l6CVHW1v61wTHRMP8BZPi2
jnCxpDluSNo3YzuM+We71TEMaFxdAy3WjfDwB7hNxYDpyusWHKJN0WCi+EfLqKofpHV5L5XX73I3
86mkr3XbJNJXpAZNGDwo95BhJAEP3w2ZInedyclLcdVnQ9vuldpKlyrt52/FzRNoqRp8AmNeECqI
P4R5ytwCfwyp+KpbsJfkcNV4bVlrMwYXbdlDQho0R32Nf6pXj26pzL+EBRILqGHOS4BIokLyqrOP
dfDqiYqcE4pXLPn33a5pWu5+oGkVXkpyfQScaBOSSUy9MbsHkECV+jM20FD8Aou2VOw0ALvptdb1
BxT4jHPc8I/quTlx9z7t65yM7lrh5HC5ErOw2FYKVSYEhkQpcJt4afODa2Lw45Osir6TIuYGcQoX
0WGhI3CKHEJg1rS35FbUfVwx2eRdDtrfB27mbmVMqC8TQ6kHEYPU2hlPuzqodOKEQgsjE69hx23x
57KlT9FWmiY9QlUGN3wIrh8TkOscrHZMNIkph/GpC7VVs7xZQMPRkTYLRdUuGrO3am4rTWtGYe/b
jVV+yoG9EWrmcz51wc8SUa5NfMGvkftU7GW5BBW7JW2Xl9vEHBT2peHqL3tAW4UIgzJcdkXpMsEM
GMOYAJVGmjIqOUlQ0bg3DdOtOegR0OVTCanG5SLnu164/o/CznQuzLLrEj+AR4ALuIDP3NDpZ8IH
lboLodgORYxPfkznxhnEUf/4TDNXPr7KhLdsUGxHSPUdNoawW7fgSrO6jH6zhiOhhrsRT3aIkmos
hb9tDFtAXVnM5rwhdlouIjsT7ZM86vqESeWpwJ3uS3qrUkjF+JLKSjv0aT67lbxNeEM5UfeIpln3
zeDt88B1ll4UvvxpGPPKMAzyItYlrJpef6Et/g74oRKRK2pag59o5sE/iLC8w90onixACEufhZ0c
so1dU2+UAsoTegLea0vFWaZJW98hHE5vVPrDbZHFVGjlMRwgAg9wr2uOoEwzNTl5sGlqRtajNiO0
jBed8zn+nK2YUQcUGZZUD1c59SQw9LxVq12kTF1WKNG5vosfgsnFDz/0ihI9qsmQ3dFZYYNORLYz
HjFATMLT8P9qGirUTu+B4V/MzDCsd+KGEJPSVgmRFN4HU1yGpvuxs7/uB0Rao8vokyorKHJgRfX8
eXkExkwTaYQ/euq71QACrl425JICdlEuWOon97XhO8wrXkREYrSjblPEBM7fcOKTndotrwKFoN4U
9DcoYBUsgPhdci9b3DaGqY3s0d4VOcNU17diddLCeFGtclQpLloq2bF34jPfBeJhNKPIkrsjU34q
mPXE/jFUev6S6xL8FE/CDIX1jvCOM2ZB3oOmqhjfN+OYqyo44umxFZ2WwzEDaEnry05Arg9gCjs1
VEayAMoi+TKPXXefxUQxyAa+a/yCDPXAdLoXB4M01fSysVEL/mET2UOMFb+ouNwmFAaHu4nfUE5h
k2y/VBbAeiEhg64ik0DCXiYqXobUTa4DYNFE3O1Z1sqyjm9xrSIEJ66dcfB2krJ/MI6Tp2yjcMjy
RQE5HNcQg1zNaANJeJJTTJQFbMhGRsf4zVOrM6i8JCJkqmpbDXx8cchVuaKkEux7/oRwJc+TwHed
UgauS+JNUUMhZtkDn31F7z2EUYDCp0Fuul73gaTPB1Vc6zhPjxQ/MZWRVpCcij0fSOAkw857+FJP
5f0W1NjawGjPoyUPXRivztTUjvpeKhRMhKGlHd73w2dt9KZDl/PiyTdVSklk5el4pEeOtwuZIPwI
2UaBd0V5fyuGSPdVbWoJaiYhtgsxF/dIrIFJy+HhhzXK6PcN39RhL9Sy+9/QzCcKycNFwQ+3iM/0
5V6cCvlbEVxM9kSjSf8X3iv8qP+7EkejTB84x35ANeC7dsm2pFMMNKE2gXBYw+41Nx0myLJLeB8G
PED6yX7DzzJbe85yU5CshY8dNZDSc8Qdeq4O6yspO4LWWCHRdoiOuHC4BezI7sQ+KLzYCxtNNBET
HfdEDB3GgiRQbRs3pcXTCwai0jpXBimJEG3XMuCfweSN4fHHgifOjK6aMCFCUzRZiX/aG5FWBYfY
3z2hQj+190+vv5oX1E4xGg2OwNc8b1F4Hln7Facp5GcCQ3ZO+VZKVoQKIw4MGh2KL4atUwEHIrsV
T0mRp3+mce27g6+cOI5amsy+noh0YoZWA6vOS1MkHP3qphZKIFBRa1U3/dDH088bhP0ODUlHJaPQ
fE0qGIKYyUM5W6TUe/PKNw765+Ev5nXdbFqFTer1pyDybXd+d0dNHcZCTuagRIxu+ZxN5+2V3yOe
yhQ5jZkFvLi1FzUF+rPWPL7x2IXCLN7X1n6gRaAmf7SKkiUabfO1oRsqaHMm2/v0+XYb9ksYJ68q
wO3NPeuQmbbG7rj7sldyXDCu6w9L/Mupk+4HDNukekP6Tdab6/P+NCeM9i2lmZ7o0JA4ztM9T6Oo
pe76p37a/1ATmTVlSlpyCiod6eX5H8qnBpr/i0F3QPm+GMoJMgFI/ANA28euLyaUQfIgLkPwanXx
5cD2O8R+uWnUFJawwiP+h72SzrTJ5Dh6Rw1UQmpoZc5yJvwqe+HAExTWjSABBgxHiO6O5XOq1tYx
OmAlbiuXjTgOh6KuAd7xx7ivo+oxGdDby3zYt1EAQ3fgkkYPPHhQ8NGJfxXUObWXtOgBcri7Hs0h
+dSnp9W0O4LOj5kzcOmu6jSgP2GmwoZBhsIQ7Ovs2MaTYOZZqzM05UBR+5NGXR9vQDX71G2xtn/9
C+QPXFTSF5wOquQwP3wDZB5mQLlnE1hGL0qbGSoVl9wfMjkMk2eiiCwQITDKUJztHztT/9qJ//qF
xc0Lj1p6yI5h6vXl7UTUvfFyO8fIXP7WOZz84qM6ZVRU12Rauh0x4jFJdhtldU3HqHrfFBz3I7fX
xKsjcnBVL4EhgvXeDCJAbqXSVCHfyTIoMVM7hJJJNSh0xZ1RFihIhsIDmG9hhWJynpBJdApa656G
V6AKfaZfEgIO7dw8WRUZD0RupDOp+zP287aELvfm0cGGBJ1RcyaphOEqFTw8+TI5k6FpfZ0B74ih
qkuFut7+J8rmUw1BAEwMQz5/IUXwKlWA8PLw8sUzKi5HJPQ1nkdySd0J/KF/+9dxco8zTelvOhhs
WR2z+PjIU2lVKzF7djtEzgC79cSU9cIDUiVqzK6HSW4L9HImZVvLk2i5Ii+L/wNcJyfYA3zCQojM
BbXRwItjolSf3n3xKyn9Qt2knqdsI8bGqEkfKtiJFx/+s3BATZa/Vg8VWlupOx71LYtnrn1x6Iqt
Ah4puudseeZRwkLDC//OwbxuMf6AZgXgAcEo2Tz1vZb4FnmbnK6JTf75z78fUnmOPs6CTTNUkTtY
I6X+knU9SuAJadW7W30Z2Y7qxfl0VThJTmshNbAOESr5Vc6Q6Bj+CyKEHzfX/9H/HHGvz49ixYIn
reTpNec3GZRNd+W2OHyyhpM1PVwihA5rxESt9tAgzsxgFA26pa52hIRLlL+B6vSgaLwXCWsJxQhc
Q4/pddqZ1KKcUJwW07kth7r75/+k+yhNSxXn2H8X5IXF9VlDAYe9J6t3MX9Ozi1MdlrUygTwzlve
Ijq6ZdySYCG9W5EJ+Jql+AujTD8euONLvReW4cmjBPa3KKWyfjQ4+uVsed8ZkC3rmIP9PaBkviTb
ZHNqvimnyB8vktAuyA5SLQsQtsAkmbzHTDleW9fva5flAp1dC1IELzi+jgNPmryiOGYP6E1yqZtq
e7OGrxtZ2wAy8vTNhMn4MF5rSfuSCD0bsq66UwgIyNw2n5s0++6ctIQJXQpM7uDG/tpkTPQdyGXr
Jekv2o7E2andBsu2YbJvdU4cRxspG8C1zkMKSoWtj5YRI7Q7vXnwrLK5heZUajVm0oFN8boJ9cb5
Rvp4XdQBoPfCeCb6vo7rl5sWpGbtQOQWOI8rhUJhrOsGOTqJpSLMpWj4hcR+yDH+vvfgnFyx6Kgk
0dVxt+vSgn5t4A4RMFNFAs3qwF5xUpPZb7lYgc86AyGodKf5Bu+Auuv5ap8yQBL89mUMesgPE6wE
VP4tTTfcde2xs/jhsD4im2zll9xCD7VyPmxWmynGjIrk2dmt2hQhAWdKGnBUauZ60iStqRGc2TWZ
rSdxkknh3GRwx0tU3rcY0WkoLi/qtZtoPBr0U48+3wW1Ftk+xiDdcz5VV/6Wcc9BmOC+5/lwzyrg
qP6x9J9GF0pLPZl4xYjbpP6xJraCB9ZKGOjHvMHqEyPiI7gkAFM3MJ0SiKvsVMBJVdI1xGehkqXB
aGOkXrVlqf3caeMzi6sqKa6876QNBSKOwyVP+qRqEaNko59fS5s2uWAtAgB5f3iHq5sVzVQMttDH
x05dcnVtqg824JMkxPdEsQq83uv+EiRjTUA6j8iZjQDFjGU1JxuJhzH12JPQGcyWRZQgj71fqgkK
/jplJ2I+8lozVRj7Mvd1m0cAkUCnaxnhWmzXK1E2aLZ2TvMH7u/I75ESiDFoBFMFYiiISyBfCaTb
Sy7DKDxoYCtl7eaxeY4BNDj8HDiPz4RVm/V2Lg7Ft79lyboDl/NaRxN+l/CveNBYXkpj7QEqnuoa
soBTuCTvYnLJRQ9DU9Oztq/CtymXLaZYsENzw+4gLS6NFc33t9Y1AUEA7PLOno/8t0kk0XeZyygD
vrPL7r6ssQ3M0c6la6ThIY0ihM7c4tuPzpaOj0v6wiS39nXxcpnjziB054fb1FpGzAiyh5GnMyyC
Hkj1yUc5vi+bwFXgAyb9pimFlnp7t0QqPYRm9+bWhT5gQtZbo5SOhGGr4vt2CNXawgevdjYh5FOr
TWVhxvQJOCYEP/lyqMGT2QX3stH6yVJ+kwliBnLIrCRFJHgY6Ngm3e7+Q2gNLGfwUmRMY9Y2mO0z
szQUqg9+ZJi4JElWA2ZnoG1nR3MtT9irfkfeF7GvYxGB86Jxy/nS+rLsVl33FEbO2y8HxVXXUf4W
spkOSJRBollDgwvMAwQE7h0w8oHfgesAGgmTYM1yhzJix7JMJPIpWeEkDVND/eHVBn00FbkUu8mt
TI1lz9Qd7GEoQZG0iPqKrHSWPdCtDpXr9OBtWbw6LNoa73R+9bTgekgYQkmbnas5pUC+CSbu5lsk
ZfnNPTCHV08eGRCUXHRl8iB9AhL2tYjc0WwXf4nKtlU6HuYV/+7lCektDkMVSvf82uXZVDP66ZXt
9LgY0NDzWrzNSqxH5Gw8ZXHfI7Kzel4FFEQ9mVqGMAVnBrB1dK/jKpW4NG4l1/cRGPsTooMhcMEy
HU9Em2C17EjSIPfL0Ri6dJH1uLH5m7JQp+EgHw4gISM4WmnSo/QrMy7Sk2LH9C1TH9caz49ZBhNj
bh6fgCgm3kL5KPMwzNrsC/M7vEt5heOWT7TdZIhy+R7tjxbpI3RA5F2QPCHv5cf3z9KO4o/rPYuh
4GaYyRAZaYz4PFwbnHzVllSMNgRmiletgcLhzawBwPA2Zox8TTiKTMbisgsEMFjfDyfIpLsIz0Cb
cqHMnmXUbBBLFPzfauK1QSXtoJGLJGiQlnnLDUMToV5LkWejC+I2aBUS6+Jfzv7zMg4iz13kws4U
q8uhJAfh8MR78cR7CB/COQ9qM81r9Ut1OTh26T6RD5m5XiIEhm7cwY1M3iXmCaghCvxHlK6J1OnK
esp334eZ6dxZ/F6R7xB8k31oQ3Fm2Fft+qoukJbAY7Jf2yC/tCIQHCncKogahB0UslZecW3Un2Ss
41HDtg7GU3G74F1Ej//wOhgRXRsShaZwsE9+YuB7WJDcDXJsmggb0VClYhLSoIc2joYDDLquie1l
pUGJBvkz4oA/A/80rQGcKq90UY3U2xe6TNQBIDtwQqDtneBPyyV7lab6dIVBjCRN7mu0q+Kp7dhj
6zCMA2I1P6mVroWzaXz/b2+4EilxFgfBAuorm5qeGydzZ8+OKWvF68gnrajpDANUn57zoTaqn6fC
T6pQvJ8JeBLxos/ewlTS5NT+Qj8Vv1hkBUdOsxlKgxj72YDxAT+V3GYJLzCeeExl4G8WmQq3SYTZ
ZArF2Ou4r21VqqMfemJHiwFTRpsEvNAtDDl04e6W8ypsBisLUU0IFw/fxlxN5ieTo6OEH5u0rPJ5
oTqcZyd4k5O3v3uwsVLbjujQhTnI4sJsJohBaP057pQgiV2eJRWH/DCHLyd30PVcth4YbphQFS9J
Xe9u5cbPHOa1XxQDM/z9PqQdb98mfoSB12+yZDAkjXHFctZHyG3x/qqO8L/xhljB119Ye0yXNgXl
ZwboBL+yFtvVLwIsd4kqoqOt6c0rA1PX+ompZyGRQVn+uuMc+hrL69N/zpFX8eajEmwnDrPurZJ4
DZI8WGst17Y/AGmbPbhN3AHG/NASQ0sv/GeSZdsaCPAwkEU/AR3IbRZ1bqsf3w2MQWzibdkmN/DD
T9K5WxwHhzW7216pHEMGpfBLQYVYGm4BxVetsjtKLwQI8lpV6vhL/4qTvUhrzJ/UD/gx8HQ26o9g
oFkb/83vNlrFRVniw9aykEMx/y/Ylnfwp6vc0Q+CtdoP66bTzarII0AMWFG4fd7cmwgW8gUzDIgO
VS2I6IxfiOTDZwJHQJJiNktkjJBJsOTr0bdhSgqjyi+gktN6n4KbiSvGlUUsueZOO/1B/KElRmWd
NzSWyW5AQmFssYyQI7uDKAdo/FdGrz3hF4SkZMuAOR0Q9cvv00AWYUC3RnhbUCVKsEFNMuCHpoo/
pEf8LTdt32PfgyqjKX/3+EiRKDhAKmTjQzTz+vPsDGatVE4CAohh6zwMbA9xbcWCIOSxn38uFT6+
lx1SB2Ww5LsdL/Tn9TtNF7f4Prh2WaO628y4uaW+CyPeJx382aO7CdN9c/x1We1kYFqiaD7ETujU
LYgasY/qMRaSZvvhK6X93tdCy6TF6J6aZegaMwmQZdu52ydG1ilCU12faTUayQIv9HWNqYaUN3fh
CXd1PS5q4unSv1YyENjsscBh8N/5BVJywf6HdjBikxsBaa5xcXKpGNSMMMtPlD5IvTyZNTTxvUDP
lKsfvBRBZKeL7Bg9H0elBgkg36ny8rAy8LVbMPWWJiJ/DL35X67lMIEG1z3mfoZiHRic/mp3wlBc
CPwAhUYc9U7t5gQ0WS9op+HrVveeJk+f+lTLBZDCBDJbDXFprL+/HsOS0jrL3WkOhZADQvL9ZSpj
nFWgcqC5IRV4O7iLYeatzlRDGZlQif2ivuX5l3Dr/frNYlB78m50RIfb9N8/Ls2f6qk2DqcvPZ7K
UNulWkPuGRLruw8pEnyvI3KhbqOx3Cb/IcbCaQJN1vsXzHzCmQubpg+7xUAGOQWeBkkfHkeVOkYv
q2UvFKAdBFLnSNLkJc9yXSwDktGiIaEF6YLfx0Onb6k4eQ4H95W6ArNQn/1HOPNdRSCAXSNSKiV3
cWhAOhK42grmyONvrsRGiZlLwT9jW32h9B64lWQK/OXuhT+Q1ooHLX4l0/mmFuU8ZQKSKpHmpAXx
3uvOPvbnjR5weJhcYxnEAhYEqJKWd5XK5tRx1ckcSyr91MlDYRonZDgKQFJpJlfcsbNQk5pkjN2l
13limVklPeGlwHPuJ2/9Br7tDt8LM+Z1681G3ryUDM/CZzCi0eobOhWRkDMx8V59YPH6T51Ogdnw
UMwVcn1de7EiFFJqAPkXAVpgDfBsMTrKgIsaVQEBnRnVQ/2YI8l3aops0aveIZCTOFyMjn9eBzwT
LiXAkzHxpNMcbyjMHEOmqA/irB/iQc17AeSBM07lfzJDJ9lJMchq2Y0CxAdqULsMBzRBh3lMPLVO
g8hOJ8OztCTgz2ZhnvvDRIpOcMJEDw+WRFRDRAztw3KvJXypzTjP4VVsKXRHKfwK5f1cs+ddlHvf
zIl6EyF2pgXST8zNyPwmQfknpVDWDH6MFQaXlBpulKlJHFgS3Tm3/ayS/SC0D7j+heMbTNJ8HI9l
Z82Cp2Ld1OGK+iueC83QR6h6hZeawi1Ypdx/joNGbwyD2RDGLzrvw9KZNiA8so8o/9kKZJxjnvHJ
jmBuGAhieahyJlgAzOE0Ro4vRcT8dlx+a7jXjM7wwubHRB5j8FfGoM+PSixBq90UDZix7EIziNXb
/+tUqi1vRiznc890TczV1kuzTLHCzzodC+cuuZSlyvfxCjgu080YoWbbACROVFERfY+NZiRL3iPV
yJff9RMZt46q2NWO0UC2vElTY1HRWqjfIQhPlgMCWQUWJMU20VUBPkfqTXjjsmXxCudbO74AZJxy
/n3dIKvEUPxgm6UcYxPiudu4hUKvAuT56bkrfbfLl0meJz1oyB2YoiBAt5P8PW/hz/GB61Q58DkB
oCLjxewtt7LT4GQRwMJ3oawM7FQyt2RZwc1ghvg6TVPSvG9ATy5GpxMB3L/oCppZzGlCR/ixx+FG
cgtm6nkKOjNhM+rZC15Soal4ejYmWiVZHPjc9CSDdranZ5VE1c2ToqgGu2p+eeef39ZNyhKl5Yry
F1PPe0SKihNdOpvtm1wXsd5dNZIs/+x+0kEf74NeSm0JUiotJFglOj0oZDO1PFgd0Uenk55JplDO
+kRITry+hC+x8oTExpRaPS6X8IvJjdCAYuwWev+tLkoqS111b5mDEjmR1LUehc2pOz+rYYQq/WnZ
N6OBTP078RRWdtmZ9TvULAYv4R4ViVdcyX8v+SN2uEQp+0FH3NPoBDqCErGC3MWuGIXU/eDAktWo
p5uzqyNNF3VV8YOKtHmC85sykBVo44PHtzyt6lVtJ4D4kp5hbEzz3De02Mixk6kYCZQhg3avrvBh
e2+sgXrQJM9me4DpzC5e6s0Rn1Z4HRGWrM56W7MGQczDW9vtFy1kSjEua58hOx36T/ZqplfI9w/F
EC40OON8VOkkmNXmrFZ4HJn/ujxmJ0rSXRWZ3hi03TcWH4Y00w5wg8JISolV3o29sas6e2/iiX2l
5n9PTzdrkIPkzV7T//YUtpWIB+wkyQmTRcO6IpDRdiw+nHE6yxLrgXydCqwBY1iMd9fVEgOcZEIL
olrYt33rGK/UmeILn8X0FIqubNUIqRN5UaBW4JvEzVDhfMhsjNeD2i61MIGZnpjjeJHlQtjK2cH8
lXYs+dd7Rnlnonp9pOJOW8LBkNwmQcs8Djq0u7oedfUOChFpf6RT6HayoN78ubOV8VhT4704ALte
Q8ywo83utL7DaowQsvDeenDwiN7khXcKyi2n7dqyC8+WqjJtr51yjUxcFD27wn/hfB2gL4ndFXdJ
kxTMMBOgHk8Aef7OCOCX5tJp4hYDadGAo20lSt3DFBTtjqCIsPoW3J8Y7QQTvEpCcGmEUKkTcLn0
pCoJ83Q5WYcM/blT5Qa/1TMfXpmvVfT4XMVXHRdMiygfu+cm8GOiUdO7zc01Wx3AMZxWROVDLGPq
UpSStS7hFEYEuingWCanZAwwVSL/frlB7XsgouY6HBf3EEaqM/MTm4pSJ8lC079XvCxxosfJNhAP
WKJR+/PNSfnKLKTEyjCL2DivOY451pqzc1d6mXw2tJWioSXvat8lp+4zVj2IjRDGYpNwba3cA8s1
Fi2HZE5b0EFgCYUiWP3iBxL+enqXfNoyOSCXFQ6+Z6lDCoXnShIiVNQJRIn8ZkCXNCll9cpoZao3
qVQbNbSHloMBhsK+OuvP0Wzb4damUdFGDTilQWpDHVBflqc7M2qByGz54n0+GcWEVABVCAxnObwb
SMUOHPktxyg2Mhlq+O2MdwHM/w7kpWnM+rr487eJpvMHkE8cnUy81eXe4yfLpajvZ/y79s4BJkY0
890uAjMtDwH9d1hgilFMb8UMoIqL5WZosRwCiNZUFvUqfea4Mwfn95gmUYoJg0f+H73giK9pzW5F
zD5By7N8zDtFrKDvI338tylmY1OBXF3s6jWvfthfAsdelHwfFxEJgrTQb4TFGnN1EubtsdqjZLTJ
oMwcBEzXXqY2wYJk0O1PlC99VbGDb5YJG3+TvK9mWt2olVjBsAkbYCL24TRrRSW9dBMbj/VTF6rm
F+n2UH6ph/pRNF6LIYhIiTaSPwi2SnvMqbsGhrOkHAlceHiUj/I1efFNKVopwAVaElopQlx2OCAt
fx6mJuxCPhZ6/A35M1gQYXHBjbrkz/UC67ylbTmxWYq8PFBzE7cv/2T4YunndWwTwAcOwJoSEJrH
j565RYHZHtwjS1SD8TeKutQPcdb1MTtBXZ9K9tKDHW+6S2fkiw9e9rEzj+qduAKgyI4hCW4oM7tV
MqHBFsgzUkc9Vpljd+UxdK7sqebUM5eU7oHwx9ampRDL8Nfz4ZexvY7e3PFPalq+Daee0TxKUwK5
X2lmVK7ip8pJhqj/ksKzbC4as5apGSd4ut2KhxC2dT0hw5DdeS11A8AFU+k7UaCWnijjW17ih3KO
44K1FKwxHrvaIcsCTvBajZIlQZcR4HXr6WHhACmqK4m7HJfNIgnTNYOTGzLsWBkBmyygsxwmH0aI
dR7LKWmOfiRXBkaNC0xDDJMoFbg+hw3hbbFFYSg8fal0wBNe9ICPTPq6Qou1KZQwL5TwjCz10S5/
tAq/IMkoJGPG+ggjDeujsXzYrJNdaiRDzWNAFqUJ4gLzecHb+aizjADmaI0E3RG13RtDkSn5AyOM
5P8wlVnEu55q/TJhx4pgRxL3aI0OEd6bLzvlz1WKTNB6vBB9yzip5maUv2bZI6pqhhAaWlsXGwe5
YqV2OzP174MPOyxAWZSXExNI4F15X9Hw8+zFIUHwucwWjJVRPGd9CtIIWa4cFFz8x5dROCEnWUuH
jTs04k67K8JP3PRYQ4UPAgVFLg6RCS3TP2X/6yQiuVTwo/CByhC64NiOeuZHay7DxX51fgvyY1ga
J7BgJHycsnir8c5NuPbF1c6bq4Pl55tfaNfuQ9/6Gi4Hhn5vWaOlYVlH2UrmsAVoUxS0oVOyRAEQ
7E8kgUMRyLKd1FDtiWHtu+Z26aJUnY7z9JHm3vvnu5+6XUkTBEul7WmBw+KNtzHkjp83FtvBAylF
Y5x2PwO3qp6Rc77LPwVjQnBZ7sUwfcaEFKDpn4RHxnt9cuf+Lrxtg9Jl0bXd7Kub48OV1nXVTRcI
IMpVWQ7D1W54ggq86dK88vr9VoF+jlFSgvJhsuP9q6OQUOXNq5aRtMQTlP9wbmXivXyB+GMeqxe9
HctKesDktWHWwYrNxvGhj5c/TYre7NezRgUY1h/cUFPr6FwLFFMmle6cv7CxocPMy+s6upowvK9F
5unUJ5YAwBLN836FJCnAppHp3zJgJtd9o4UYKH4lxsGtXlNDHvpM5H3+rmh718oMWmlpCNT8fUPt
IBddhniPA3yrjJgL3z9JCNAJ7SreyUd3K0uyPmO8U3L36wzLOPOXoKU1A8uPISf8zMVXp8xNBpYV
oE2v+r9BrMuHDBYt8hkj7YKXePz7IuLEsTC1DL4I+3bNdZ9chfpJibMFfzpZsBTzsYf7qp6Sw6ZW
8FYVrsl6wZ1VADd6sAlQwpaSyOCpXHwCu3keE56kyddU7rc37lqFgG3mF9Pd2X9K9EofG5QEQafr
ELUNPnX3BxOIpuIcNSA4OpQqqPHtzTXIzuXGheU7NGeGr78aZTSY66fo0RaEEDg8t8lubK8Vaxrh
0KCF4CHuU+C9I9rUmJhZARYWRc2GuNpZt5K1k3c58rJaFQENr2r2glre8l7MGVffV2nC0J72uARQ
/kmXggCvm3wX1wLw8dNPVj5dq+7d2zkdVBpru2wfsaJFBiAPTM+vK8mbhn2we+kBI2AwMVNA/n1K
tFG++L5snHLpJpJ7K0Jy6RvRwQFfrxTnWipuz9WoTO9mQDL+bQ/IM6m4OAKdglODIg0KI5X1ha5A
wiMJQ567Aes2VIK0OGfe1qSh/xCfDmyovL940RRTtTeW8mxEM9muaA7qAtRZeVcE2XQhDkgBU7Id
vXCMGFTQGyEmBwek9m7/8o/uVFCOByK4CzcdEvBWuOPwNyp476kyuqLtTBd/xAvi4INBd4xqvSB9
WLjz7/olwnQ9qQur9VcmrmaFBq+2BFAKD+lsDyVEmBkeBKecaRf59yZdIFCzZkxEcBg2/36WdFT/
5MbDzXjx2oNJqnw0S6KLiHhHK52uD/VTu8de++XpQRCapuRdJ/0syKjZVyw6J46SaJRhly78FzzF
NXofKNuclloSvJh+0EL6AwwJfxKcCHh/VqPu4C35CwwfmsLIfZUOTr0d/yHSGua/2qZqyLNBolWM
mGrq5K7QdIFtkDPNlvBhXatPdbdwuf0D0gINnF5XaXfRFJFAEshFNQSa9MTFPmtc5gVYbMtuTLe3
Z/E6PsTI9zpJoSyIs9/L0pgtwUYisgnCAS9JDvedmBlJsrJRKjzhiVBoCMpC7Df1MHEcC+oYfEkY
+azuc/qKaLmdg5YxdzSXcu+9hA/YnJbP2c38IrNNN5p8BhrSbB+iTDy/Y3ZOVCZUrCwzh/WxU0Zx
6Od1GvR7ZglxOulR71hI+apuXz28vZ7vq38JmNuWpXJ27k8EWCKE8r3qKFRlw5RAdyU87W5CS4ns
HzLwdRQPlFdNuez3Wk8hqSdiIH48LqE+jwnB/YQhFDXOZv1k0CufDi3s2iWceUkz4UPIQ6NAlQ3C
ZPLRC8ROHlXRsjhLrUFa4yXFUFidFIGs614zYZOkgEol3ikjC46K6Z/F35OnpY7pYWIdFCmsx0sG
Djt1VxD/ZcBCXGb1uAVtPwmBgM9Nz6vdnJDlp20HjbVknhRLGVwPtXztN3L9wCJJEgmceUOpAkP2
dW/F6NkCBeacheH1zEvavEH4wKHyDklqxw+WSkE0eArLXXbNccXdBN11j4PtsK+CcQCCFc4uXaZZ
pVHqv6uPhBtaLZLRMqxS8Rh/NJIORFr/WwpbNLKu6FgSNjZ+5/xzo3izTKs+iQ4IMmAeBcnf7meR
m5ShnrfSOEqIEijl4iy2m5Rsi7QHQAJBVoK/JVhaUmDP1CHMecRwl3qlyvqhNUfihiA3Ap2Rd/G3
+s9H9r3gZKnyMPFKpz6VPZgNDZejNZhoGnVECpvhk202j10GZ/s6TrqrSTFx3e43PA6xyNsxrE4C
RqtfDQPlG5Q0ulHawGCmo30ro+OWL9R6Zgyai6lyRtM6KonSaD69qJV72H2Lw66yK1W7Oq/WuHyB
O/ZSExNn4YL23X1JSP30xLapTtv7uNE1CUhwinO6LzklngV0WpbOZr0T4IiZYN7Lh1yaV1SAlGkL
Fjk+i9x3blfqOL30ETNSMsdEkK8eR/FRf7T9FTNdb0tjho7POcBTkyziAZnHQvNQ8hAcE7FLv7Cs
wA4FUf4OfthwE5NiBGnrUgDfmiU0ckbPjMorXqu8iFNm03iED0KRFGJWgyEjWCUIl18ihj2tKFox
efqQnOJPqj60rx9Rt9oMKMVPvg3PDJoEMshPHW3ha2lfAFceBQMWGVnpQJ6IyZSb9/CxaTQcZRQC
hRmGhCGxvTt3HnpinU1cQHFrDS9bBaBkHACnVlJs5b4p0QGB7wuFiN49CGSdDmODVDlOrLlH1ipa
Pw/OAXnHaL2RTnvplpkCvhvii/SJUsqfwgNM7DbSVz7MfrE0QXdX4nu0XhCZx9iCuyBgiSm+3+0F
rr9HbrvU2JBnt2N89+h+C1URHUvLK0fU4w2oreMt1H/aM2qQiBE9lqXKy8aXMLE0rNHULZtgzhkp
9Eh2hGQBuntI0oFhdShKAm2AN4pz/dguGhscgNCwdBqnNlKX6pa8HvRpNrOyCNoExs94Osipe7bB
LFg/rz4MrTcUETETf0o3ki9uuUqF7knZLKPuNznjqbwYxZQltoqhFsj5+KqMVVXC0wTsaU4e6EPw
1FcJ5bgxoJsMpBeKt90j9NVRGu0cz0ymMfutWY/a0rqLLaqd8bOe35a0CA/eDVF6TFQmRgIpq5k7
AnpBbOmUXpYvnSW2OPIRdu2DxGa1b5fvom2ga9j20ClJZqyzsQrnx8tDx/TKHY8KhLgZX10s0M7w
bEo7hENyDMvf4skmriF5kSus9OQujEM6gDC8HyRldD8nqYv8rFbU9vPh+7J4oLYYTDoPIlwfVoz0
8uwtL26JZo5YcVATGPeU/vTTeDAPcQTYmQyWXOPfxyMozoJnAtfoF8b8k90erLPg6m3dGrag+Bj2
dM0mOzApB2UCEz7LbqU9DDVLc1AGJZNQrJ8Su0r+8IVTDzAVjc05UgcsKyA9Y4jbIAxXYp8FCX7V
/6eVNXpUsc4sxHzI9ZL0dg/35zkGRia5OHVYMSPNUClVh2lWB4yPzygCxgKT06idi05FLfAyuXfU
wILbOqKXWNStl1qLKRLKYpiKD2ACq3tucl+iTDpx9C9iDBV0xJEX+K+BWcm1OgbFxwkXgnk649XL
XTgIT3MC76sNcVHBvG2ijrBS8j6yZc7XAs+1wQKoBtL0Y6zSBB0FbxK2KS8/X05md4FZq8D33tce
ht0/1nUwaRkgRFtu9J2rGmNtul/Jo6ZwR37l4KJDobWFHW4wa8GL1ZfOePHtmrmAbnhDz5mGAR5R
dgpdypOOzqGFVlwhGZb1RP+xvLYcGJV+vKd2U5Q8nX+0FHH4bq/42z+rDpNRxU5yKpn2gGlN0Hbt
o86nXt6BHt+AgDKw7BCYJfUQ0u+a2g3kxuKV2fvFRSDQgEv3TNTAIOEJF8h0lkkT62YiDqArYzjH
G97Nv7ViJm1GgGUldfPGc9Sp4TXZhjoAPswrV+JOziCdoCvLlp/9s7H84uU80Dz/Xai4gnHe6mWM
JQ/piCPnnreF/AOCPnuvPJN1n1JCd7cBXAUnfbOUiZLII/BJohiuHuUHvgPoooxPrLi3QN0j6WdU
gUvvJY72vIvo/QhPspc1fTAvb3s+oA2CiJyKiVP2CjDS2QypeIP90OF1z5ec8K9+ap4sZKp8SLr4
qVl8ej3pNUI+WPrKG++Yhf6UpGcAdSM04WxwHrxol9yNqF/dwlPNhmBWlYL8Wv761nJKGQQTxc+F
sLell/MB3WC2pf0xjs6bZkYsbnQ3RShDwRmj6YCVktln5s0s0mIRBldiDjNSqXl9QhWv+bKHc/FV
t7Uxq24mM5MjriSZANreAdoY+Qq7bqPiDmPXRtPeTgbTBONlZXVT5Pgbp5Rw4TWksWDFm5YpNLc6
dwhiSoGZjbF8NER/APH6UlSJu1DE02NJG7ekNEYGXMDocXynIkHTXHVvnzHeXKX0WSXrm5ARL9l2
w4m7ZSE2Tz3dT8uL4WtjsLSNl+D+k8q0yViYHRzqRJ9CSj9qQewug2hla/0vaBoommTlxnaxCzqK
NEVwGRyZmT0goQAB+lD9j6kwpnENf1dgvtnQT4fI5oRRN1xLceiR+v2pikA0QiSk1vE/LsMXpal4
gJzUPLFQu78l9l2d9XuskaHYQOiuzBmUKCD0AQL88n6XFxso9zOxOJVYFDyS/xrss75ONBgG+8SU
ZvjojpLgcxD1MgNGjGxzYEqbUUo9HIjnIdcEuFDBtTTU2sqLQvEJTmbA2lbn7st0LmsjtwYplCWS
dhKufwOFmvq4ACJyswVI1OyNbDTczadHC7brBN3S51KsnMeCRDqEzUZuciAlwbT/2RJ6bKAwBbFd
KBmikfULpDDE2aWg7a0ScUp6MoRGcg2DRABLODK0wo9W2BXlKnKvLMhk19pVWdhgUBKO2bjNx0Ei
CIufrFWVQ36kpKZfFjdZsUz225/vWX14HMsLIMVcXCrXwZMnCoAmRDLbp7Fe2nh5dzwHCeSTPKMl
6ZvpGnFVXdiZPPEpRUhbJM0MwugS1jpTA1gUpyPtXQXDdW8Teit8pA8M5OmxmOR2zJ52QtBgTwSQ
KzQeT9zaZDGTiM5MF6cdfGNm1Xwt9zfaoeZ0KIM4d6NuTN765QLzyeDKk74nP1moKEuovEE87HGJ
kWZs3F9Azv7wPNE7+/uc6pm/enExg+I37rCLd2TLheO6NSCdxFOvweWg1Jn2hC/BtoDbhceyT7u3
CeXKZ/CrLY4L9N9DdDUKlFZm4viZChaqlLbzH+KFSQGUS289z+a0qexcwMPdvpqIiNETHbZ2z/IU
PwkEb5RPRbM+KiSrAmVPNBK6EmwvpYYVdnb+A7OLdlKeDKVZruYQ0/karkxNph9AE+fh+R/Y80LH
c6ZSroXZSixNiS8kc19J4++eERu/g39cXB1bdF5cCSc58oeFQJdsNVVUjxPMIqRn/3yIoG4/hl/P
zu8wb6lQjOQ2jjimsth9p23inqyB0AvZU4jR/emuLmyNkI0xEjVjU3weezwjYMTaDEyIaYoL9sL9
4n0s4sOXdQInItoJygI5G9TWlHy3LGOkdrOlzIGUUiGDC75Y/XaKFqbBa7C7eORUA8DFUDgcDrCj
6EfnTl68GV9pik9I5USacSZVf7myS6ETjo9Z8H8OIzKF0c/goH4wQg2gEMMuM/MwwOEuEPzRBKRc
Zn1mZMeoXVGwCwcm+BPg/tM+zDp4bqolIsArarB232pp8nR7mKgROajNyF5XTOfLspY1mXY6gFZX
SrF1ypqufk7Z4c7hPjz6nahUnUJxpyd6xZ6PSZT0DnJNVuOqOYDvChhfJhwAlUX/MvZ+T8+wxmZh
YdU66tQi0kXcnwJq4O+BLn9H60Infh2VcjN9Z9qxh/yI3KoGYFsUEl7zu1TNkaJW80ItmVFUDtFu
Mq0nW6HXd65FSdZj9RGLkp053bmgi0ONILckQTI9xL3ryfJj18IYUGNUG27XzzdxU9P9a5Ibh4qh
OpviBCDJ/QoO+JXjzQnS+KAUK6WXbB5Mf6rw0Yq0hBKtaBP+gJT/v20xwopA29DACtV20N86buIJ
DUdFQt5Sfocj/p099IMTstaK9h3BnV1qrEQ+nxT7NoP4T0v6NmjWNBFPe2cLdBRpElwO+nd88wVG
AGh1m1iSZB7MgyeTbWCpa/T6Iyl4CyJSN3BtsL6egnaauXjTD4lYTpXLwp7qtJUMZya+NP/gGWf9
mZA1OCHn8j6cWZ8+xoLnhLV+mvnAsBHcyseHzP3f8d4ueV9VsaU95drH1wwj7/v83KkIL97idth4
NnMSPh2aUwlxzg5nRFjcnEECo/jS4AhSQPP6HCa004v7zg+duUMbgZsS+vBFLO0ZDmt6LVc6lAiL
8qBRYO90meP5M508H13A5QqQAMBwCINTB7xCKt7ZkEsyJdykYHhDZwsdB02TQvT7dmI8TLd1/IZ2
LnNmV38r4CHC3Lp6sv87NjIh4IwYPj8SPJpQFJr5GQLoFeOuIJGyh0fd9TmiBFCjE5QaO9kfVRRT
2zx9p9VlMVWuSfINax/L4yT5ZMW+Hyzv1RuRxuFT2q/jbnq5ujg3Q6GVOK4J0kK0Ldr4HvStER0a
ck7LESx/Ziy+26TRLqiRH+I2N9wTPcAuVTFIrIxSTYNM10+tIzcRxtV8YHIqP2cKM10Bty85+lnV
iGLk+UzPrcbqhFN2RYXR5aWw7VDt072rURhrgliMN3FruBKDaPXC+8Dkzinp+UjQvDJlg7TnjiDM
+/nNRFGe+AgPY8KHT3ackx8mPX6SDGujPVJSG51uFkOaGifyOtne7zpv5ouYiG1CGSLdZrNlaFAl
mH2jA/Zy1CGhsasKyIw5Db22BtOsidUBePhVqH4w65b5tGFHBVjzNvdwnt7fyF5q4awyUQiq3Lp5
UuQXdJGKcc0PkailvpYjvXM4/LyYf1H5AhHiIRDMcMhdujQCRKPHWQAVvSJb1xJ2YgI/dZ9fgx78
do1+4Hj0fGbnQlnt+5pd+4mWq9BvsM22r+wiQ+L3cxaCohuubtjDTQFmihohJwx33rNpNWMQ54Y0
+Ez8gWPslQRj/fLO4YCZHpsLd04GzvtJa1GKuqbBfL5qoVHQLITeyLWUlXspvalzyKVopnBDz8S9
lh1W06W5dtLgjKOdyGQ0PDOIbGL8fUtKOQjsRGREgHmRda6A+yPOBkgzHOtR/5yMzfQGLL5V1gt4
YhUFGc3MZITRKGmxrqyE64/EddJaZdhJkNZOntywxC9CpKv8GmSB4a5jM316u7/4/ht/bM7Ath13
iMiaOAR+47SVHkvF3dipARwpj06dubT7vRMtyk/yBtj7gHwPlzn0+bSRQLJoga/NyDbD8mT6ajs5
R16l113fR+/tBAMZdUQ78K/j8YkcG0PyzlF/iYRRE452NlhNAH05JDgTE23q32AN7FO1zLkWCY4c
4iD4zC54uYk+EkYqnAJJI/kxO1/jBgO/FgONuTyusw8p+OM9/XkyudvUVx6iMamE4On/kk0szHg7
p2pyWMIbZ4vsYhaL8amXA55ceJm2reKgDx7zrs9wkW5FeSIG5/CmmBR386gUEkfj/7krOeywL3Sj
RgKD6ljuSMZ3BSx9GMwZLvxzwNwD6b6ZuuI6fQvD00RVj8q8W1P65Gx95cDhtSuvR8XUexjqxhl/
PfhBGyYB4U9I7H4BGkENZc4WRL6UlOb4y23aZ7wfj9t1A7AJBMnIwOtOiVjAFCM7i3zFajLS0Ry0
kOLPb1Z5qUo2Idu2HLjqMfcMUNCzV7ANtrJuBQMyXs6MQ/d96hxiW1IYz3uFo5/WYOhHRm1qiOFO
PjDO3av1iqCcWGgck67hU6qau4jvbIoZkjHji6o/c/S5Id+/wi4Y3055YsgkA/KX+7Pl0H/3D14d
r+6dqzsZJhALbHASgIcwyE1DDW4wKfHOw6/VID1WaLly3Cn4uYnX7Rdm72aLMZtJlplSOZs/CXlN
9/TVi4DqwHDv36JMstvyfYWV2SLCf9F19gUUxE0xPLBXgvtv1/vD8UQuww7MPJrExhUEHGJlu3wA
YGl3CI6pwhNOtySl5Y4IDdf3BtoVHNzLy8f90/q6T9DIyaNWdMqYmESFOVVH519ydhfcD5WwUtn1
ugl/nCjIUUlrrl81YcgouLAkbd/+o5hEeaAJeo6gV8TPFDdf2UyjTlA9k8nP/3CURprzaH8AY2YF
cF1Fjpb/+fcU9HtgjTr4NePEyx+HPYHVSkd+Yv1kJJJyfg7GnarL+sigfrt6yIiBwmjWVEV1pfWn
j2hdVRGJkAN80iXW/z9LhHCDDcdJ4outeJvv0p5NCjYDQoyhbvoQCfezwpVXNJfdjFERqmd/6f7M
wjQbes6/Co3TkOizRUDlGBEQENkMm6NJCXlFu55vdOmQrk10/Ym5mIkVJUOqUMI/AZAvuAT3IdR7
hfEi1RjY346AqN1jaRFode2ypX0o2mmqEUIQCmU7OPvIxPyDhCS4QxqSj+7f25nXFPUiSOzB7vIR
CmiNP3koT0Xav//oPabZYF1yoQ3qCjRE70e4OzCp5AVrWEjzeHGPIhHQuKMfMkSZ7xmMiu0SrEhQ
N0oonnS98GuW44gUAvejTiQyiPfD+TNtpEG/hf8JLc7Y4TY5khpbbo3awzIQrNBPqSn0EtkjgFyQ
COy4e21p98+2mO0z4kivyG6SgHM+a1SqLEAD0T2uDw+w8BffBQvos992k4jc2+uZrqJ3lirwO3LG
MxpCsoewNokbJz71y2VVc9OYi8q8a8e0LQE509JnlBbZxhI71MyBTpJ/3YQCeHtHBJb+StZ/WZnh
7dlOhjXPeC5CxOml24/d8ygnrMlg0ZI43V+I14TuEIRRRS6w36YjnJfSoZxaJ9Www6SnMMbC5tg3
16BWoWxQ8cXkxurOH1wT1e8kqeVgVUIik0cf5p/x7YcqjM2mXP3hv5SwPRPRf9juvsaTRpHp9hZZ
1tHQQeT4RUvEAVJ4nxtRBCAGVTskfbDmBdAnTXu673RemhodNVXxUReVBRyRxlyl9jPZph4aCZhX
O3H43XEcJgVrfQmHxYwUGllJD6N8OEb4VBEpF1WTHuOeYEcqHg84pHq5MWix0VP+5PVVpQ1MUnLx
w5cvAys/ZJ+4Jq7AEeRVRVd5RTCCRlJ5ywH4xwMvXbbaB1AegO9d8vXQmOhZ5kogFKQ9vrkg5ke5
QVk467vU+QN9y+M0vwydBRdrCWbaBUh42skwO3YLHXklL1InU2Z640twOT8TF6drhoUZuQ1nJJBW
jhuqkpHP1kmEYp5yHIPsxxFbWx+aVHHcy0KWIrk/ks+iasRZ3thtnUc9D5DilAzDFdprJ22EtiVM
no4RrRtLHmjZ2HHwFHHMSqxxeqb2GPhJhNunq+7mTveZetViQjtGo7FdsASOHJrhIySK5/3ktd8Q
dk5HIMDVqoPc2GcoTBWC4bWWsEtJCdRrsc6mFHoKBv4KEpt0eE0TlEJFYnd7JKb6dMZxSsr0fFY6
Pf1wUi6g4Mkt5FVMQ2w8ZS72shoqXX/6MB0O6VOaMS/sBLuRUjj1OXbnFeno6Xt2ij3vGE9sTOdW
iwx4Q+gk9or/L6gdSfP7Nv5AWknU7iOSEeAC0kkxWDG9mz63kIjeBj7krJ40/xUzqc/yKuSM+3fI
lO9AnJhz9FvOPVdGbwGwNfwfdbWUQadYFxwbtvBN+r/nGRJH0U+lp2DfqWpMaz0FBuzxTMd51K/0
Z4WG8qlOzZjrx+Ee6oqd1i/hALNm53PwrNGxh9e0xHjDSj/Z6/TtGWH8VVe6LrpqJ3/8lgmzONoJ
VxX3ANLzg0Jh5HIroRHMGL5NfAEBd0pKY8R/uVmeOR3o1D2w6tXP3JP6flx/yG/Cd6gP//xkOw2v
+Rh4iJZjSpRc8iHlSXJbzKOzWPCwojl13QiGBJRxRvJN1S+J6zNW9Q6DDAYiTRseXhF2w3R/6+t4
J48MXziuRhJ4jOUDjlR1k5teqF3Fmpptq0RSl1ZmlNjlWKwsM0G5Uu/eGShJTNNqf6RoecdWiCrK
7Iq11ZIe1REwz6VwcjbfETR0wixBlGdf7HEXAVzjmSpegGtWJ8h+9DnOSJs8fSuTFIJobPuIN1U5
soksphaXHHF5Hj0Mb/S90LvGxVr+sut0SHpunlJ1ertmMKxAM6eagefv5DS3C1mAZjdfbixg0xkX
aZ7BVqEiWit2JwXjFLktmaTwyyN43LzzyolJOFUFgP8v7M9MGF4KNx4kqzp1Lh9gsVVqTKC5K+iQ
YPY06qYMChIKvEU2+TfG9a7RxvArwlI42y3zwMsfCLYBFpRdUFGzUIsQ2H+eIJL2DYABbHdU1yb3
W+gHqg660bsJBIOYHtNyKOHhoc3n1b6c+ZnrKnkfMthWKuFMLxYfXaaOL2MOQUIETQw3X7kefiK7
tdRzlC0mzsg9g5bIbzAIkX2fGXWvedN+LJpaGyIfjA0Y1M1JJfX8CEsWJh9roisRqKoBW+bL0Wnd
3eFncpY9EBg445f3BX9u1o8NNgYtvzZML1qxnocmYQ+QKCgGrvYZrf1+q+LmT8epb7UUSTG0+rrh
grLRcAGQ9vImedxCz17u/Xovt92iFK3OSJN2DQPd+swbN5M4JB/QRDTxRd1svAjjbEtX8BFN9lCZ
z7hhzpC3X+MJoAAcObCGDA4JWKfsnScjtN7ovuzJ25Qsm2i4vt0YzUcoVTgwsgPud5dOENNLhCAd
4hPEvUY1XDb8ohPtJxQBFgTD9OJS3ucG/UXvwJAdLJl+8zxSZY/wEpX3ckG5e4Y+es2AksjtDMC5
8EjBj1gjl7UESdsNko23BlDXDe0XbrKxoJwIgmclZx9igZp7DB2JjXo7mI1D0Q8DPwT2lDa4bzaB
GFN3mHiwnW1evSUOQ2WRVJ4ZlUqWlSKxnp1Xodnm6wYdgrXJbWYb5hc/dugIdmRCFwFkDjX5rrTv
Fp/fjz9QP46ym2arhNvbvthRaa+J8fSoYaK16AYjXFZb3Q1iF4YwCbqEnaGQKNz1tzoAhWXTFqQr
iSA/0cQnRwLTJ6okryNu4AsSKOtoBJzLkBxyuR1isigmi44N7i2yXhZPHTtjC7QKTuXAiXRcywav
7qMtSi+9MSa0d5fy4njO1otjZqGhuV/B8s3RLI7sVWNEQ5q4uEqstMhRFPR2+Urcs1OxzJOVW+Wt
t/S461G7bsPsJYyNY84+fqm4cfB5THDpXh6xa+aLA/Y5fFkTPs3vqFezP91WfSgCddrFhinPipnV
nA/SPJLMvIdp4CgsNAvZmUiHbBoO30Ar8mz9AZpEsgHNzTFvLIMgzKpQ5oLxaBfjh42VaGb8IVgT
6cp7APBA01B6iVqyWXgqEJQpC/Yx6cPj7ehmVn0TPw1+T+OVZp9kQPYtFY0KtKuTsyjalF9xoFSS
edFyoJ9GqNgG4Pih8Mo0KIEh87ZM6Limj88eyLPkS7wxZHwC84qJhYvVZw5/g4ztX5rFVo1x5ado
xzpWRJocfbB1RaJB7hh34QNxuwgyCswsoBBEUJp+eUE9jPXcLozZ3U29Rjg3FEhQml9G4zApmbK3
9AG6ZiUHLodqFKq0KQ0ExyyjVax0hAMC4L8hHFddy9DMqLB/rwTHBYkeD2jDfMPijPorwjx2y5Ve
CIWlX5fnDnpJwuFNZCukTpoSt6Dc0pveifV7cIT8UrEh06+wVgMNAchoo0DF8yNtjJgeNNIAIzkG
0bhnW2xGSAC4PP9IFfFjRaudAZ3bxbcvNhoSY6rVWws5Wu2j6FI/WXxU04qykpOTphkmE6Sr2hXU
EnffuYcp5TsD5LIcx6K9595GetCPP9PRQ67RDCzGqkTiQgltzmiCWV537COsJul95E4DJuzSWsvM
zt7kVX3+pDiNaXfItsCWjpxe1YkkT+yca2Hgrh/4KlE1VWWD5P/5K4CiNV71pPRv14bCMj+4jbkI
qiJ7HvyVJLL6sqFbyEsQ+UlK3cM0klETYqmpFuxHlXQP6V9DmAwH25qWqT0W04VYysrYoIIKTaIG
gCHUI0rFHxETqfwYdlC3/SCuMckhryKH6p496NL2ypO16xVNLAZqRCIKwXObksfptnOTWhv7Zcau
7/nIbtIYKM/qNXWIIwDFiSlr3fWnmqm8Gaqik1jLl4vjtEepQwvM9MwhKh9wlErB7nht/BBE/qFN
6EvoNof/3sicZKEt131HPpsmZ7uxwq3+BXx1cquytn5bnYnAgidE4BL8YXfXOS9oN7KV8RQkCmSh
FV6cuYaZaum6IjQZgWyLT/6uFhGrGrv4qksrHOc5BRqKJJgCuM1A9WyyKqX9pTiSTQpeanuPWR5p
EuWJ2ub4iSPwzHVMnn8NjBLo0WFCXuAM1W7KOiJ7uK0P78N24Sfahh4vA487NDeKrkKAoAPVoW0r
TOnIUk7x+q01a09lkYRciDSQK3HDkGvxQS8hPCWvSQfDazRtNLQwVcSlP16BZGgN7PkDxwYO02fA
P4gJer8+4pS1uAZDfxFFy3NQPynw7219XNz97Gjc5KY1NmU+WZxQhDa+RfJWHgV9FBqGIxFjADrg
/P/5QoR6UwGez5SeviSQc8UHfGP9r+jIh3dwR/Bc79D5PO2CvW67vMc3hy724Q/04sD24jS3pbvZ
M/89dmL8YEneIBxvPRVL6XsHcaTOHwpwQpFqpdDfZdZQOYgT89nXVcquvLpFDdMdFAoDsI+2Ikk2
459A6DUcPI4ik/lxv16pk2gBQi74YfKAc0FAFkS7+7Ig60MooWY+6357hDjFBb6L9de6C3KVZTrG
rfR+uocefK5OFdc+FIGWjaOcnGEnyLIs8Sv836afO53G8vmZqFMbsLWGLpF1MQ47RUYET3HVZaoi
e1paSEnfbhBt/TPFTRTMmBQW3cpr/y/G1VM8YLf/ZA5gGUtXcobLZNifnrXHHx5yGRc7PcTZ56YU
r9j1ghOEYFKTWhsyiLH7Uc4588gb2uUR1lV3+wKgL5rnsXQ8m2UCZMB2Vyg+S6rotHqxxE1PpSLd
HgozERC/TRdt/OiRUbh9LHH6jp8ElSscJV/S5upYw4AgtqQRMoz0+uTGhNjKb5ZbPt/t4w95dMxl
e1W5gfD9uoG1kSdzfXeFwtF6hc+XQtxI8/1aPIY7qfiFgHzV4peQeKwmRKC3wbGRZFbCsJoRo8Qs
wXA2PQcgMPXW8lPsTa7dBXCmUHi0pvt3jM2Ql8ayIuHmSrF5UNIa/k4VKOiNhIfnUSrv20f3/JIp
S+BzrSFfVsFjoSxzeX6tp/+FDrvACYjMTcrUxAYfI5onCxy2AvQ4kmLi/BItEuQkSlwDS9hZyTPL
u8m13LEGEgXNUpEwGZpXrGveuAgKdnZg2Kg2LhgLt2kIcQTDOn9Ds8YU1wzwW99FpelYlXPM7aiH
oSKQ+c+IHB1RD0Lg8Jem+/ZBJNmDtleR5Xj9tzQm7WsirSqLyygmUrSVRu0541LgkZJnk5p8NO82
b3Rd5vllRi33OqLGPWnUbTKD+g9n9iZgKjuh2m1McMT1jXfal7YMKulXmwuEel+guQC18hFGZcbF
EqdZlNcsI+BHgR6RenEx6xd+0ft7PxR93kQhbBkS3M35QFldyCU9EhD73yT3jTWn7+a8fywimSxm
hhVhMKN1sa1D1Fwci18hcZcplL1MvQlMyAL7LnnQfZkEcvyIwxa/14PkwO8ZKeN16UVt3GIjVov2
Zy+mAt6I0/eMqjb9kz4iGhEwpSym6kek7f4TzJD6Lm3+ibmhZ9XU/DTzR6K7vsMqrsAXl+ZaosNN
vicfB8U97EBaOMbxvoz3g2/wBboube9itnIGifPOtToQMrGURSe7qZ5Sabj3JMIhB0Q4IFaSOKym
bs2fWEyklRJBXLIVTtd/9KdhsVOYQlFkQuJtqHTKUZ0Nr0NsCnLF3ffuz6NgWrlP4kUqSy/SIa75
m3m0lI/w2Bj+BZEwo9I3RrxFPihH8eQuiM7j5s7t1SxbvhcRKlVbUAAR8iyhDgBRAn4a54zTk1RW
kZQ1Of5lVKO2CuUaAtB9viV6+mZw6Kgqqc+wRe9QR6OI094vonyDaZYOOI5yLvwqAAgPlIZcyfmk
oyBEZ2YblOfMJ1+cfH+Rq9ZWOnmVpknobZmYAkFcTr7BrmYfGjDO4ChFNgZM8FJ5iB9yIIwPakVV
EUvLgEiCWIGiKcVaKR1lqa8Wos6NDhzqoMPVP5OToouFy3tss434pGOFGfKaJYJxirf1PNd82664
aEgoKdeoJw1Klorc6xHjMinVPS54qP3CEdab92DUsF4esSLs5NMssyyjEmPJjaIyDJ0HPWLq5UvT
DPUT8P91pEoGGOw3k1WYXvqK/Z/gC6JqOqcwLgL5UIdh1iHI177m/D+01IIsf6Pm2piohDgjb0rW
LnmuMXfQlawiXO2LwSsN+86b146c6YFFLGLIxXGwf6RKqhIXq9ckhDs6aqp9bWbIBOX2Wb5hAtqu
KIrAzjRWVlt+P7Snn3EWyVIKxUvGu4Q/fC5xTGbVjq1GF4UXBY5Ie/Z2ecpia8LwPZ/S2my6z8G1
QWq/4/+wPeQLEQ+q2SzA3EzNivnt5wxIohYnSRqkY7V7bAY4htDiH0tpdTP1FQonLXZ8j9OL/7p4
zkNvskzNfOCGp/myRVH6e+IC0weINJlJ7bAAm5SURrrtS6gpbKX9VwWevfNNIapRaimValEkzmnA
c/CiUz80RWKCAErwabed1t7tdFrCV5YbQWMTCwY2MEAQD9GlqsXCeYIG4MDbedN0GLU9xq5cH0Tc
bFVR2RVHTeuBAmOSzJnItVWarKg8o2ln9Z/Zi0EqPmc9ekxrm8vNQq6Ba/C0Aw6fZWm8uHNcmBAT
nDYx86rFX+ZUnjtFQukMbTA1oaKgM8mcvPKytX3738D+7U0bA9qvB/V8Mh6rVPVm3uIi62HfrTl4
8g0oyJx8A+ow0eGhCPKtJl0tjV58tCASClh/jhpWBI8001Rveuo4vb3tMbIn6LQqKlO/pLMQ2QpQ
djfgJAaMcIrIq/uV0psx8Ln/2AjNcaF/PrNqzq5Kgpc3mFrNveWeLOFAlV9Dusr/ny2qmZ0w9v/D
WDta4xsNZT6O9grYyZpTOL+jA8jaWOiiEhtQIfsrv6HSuUa3tS/ZR/Xxg2sOWywwhZaWwmjn+CYc
l3bvk1peS9vvXKv9563hTyT5GCaatMCzQcE11ESiIGjjPKfFllYPyktdS5g2xKfCkQKZHi2zQ6Z/
dZQLlALu5vXfc3NoCtP3FXNaalgsu/C0hxPFRwBbqKnCVT0/d1L2rZGzkf1GsBzExuuRaiM7o7b/
s9dEJTv1RBK/td8UKZgs5OIEkaGwn7eQfheB7fv1vqoFSmRMHzYOe5/2uE4XvK5dFfiVopCpKNfc
4uFrrHxqUsjcfIbW2T3S6g2P2XkaKN6oWwH9B1bPYtjVd4VrpDW+dtTkAoQEIWFQmCV/9WRQg3kT
mW0OyUp4V+3M0Pc/+tfTILThcPivdKyEKY5zCv7wahZlaIoNZXYTanK2c/YDNZcBTkL+MXE8qgGt
2XGslPn7aCwT8ounb22cjdJgEfP22E1sLEDZKZc0dJYVs0OccKWSAjTbUueiehIO33xJPK6xlFLL
ZdYE+jp6e6bwYpuK5D6xRryRrIylSp8HNyY8Sa+x+ej4L+Icdg/iVwIbxrPT73N2otxffX6FKbkD
5awSd7uEouPvGQ3kUdgfXiCNWN2nFDL/NgeJ20Jdf5OQvv2RofhkhTldWHpHHxRo2iDh4PeETAPg
WvbL9Mu7//y6c3fCWLDZsqoM4SLUlIUruyoaBxmLYaOCv48ZnrSKrx41KjZJvuqmcveDpPjtZs3f
n8Pq/KSCzrGWzadK3ftUmjS73gqC8BRSD8H+wBwywar0xFIr28eQi3JdnAKYul7AhqvKay7HPPnG
W7LpkjvILme9EJqSGyf0jWkkFNljsYYxoc9pWb7KuOSNQl0cRy4G2ODvRjKsiSrHBt0Z1a8+6xTk
Xv0MbH6e4+lJgdqtiygFkXK7Jdp/F9Ll5Qi9LWmKyQXA6G08iJO2MUMlSU8WaC+qTGNupZPQtFdl
1VeRjDSpl+uwMsicCpRUc2oe8t/7MUHoz8zhOsw5E4v7kYFUKEVVvv4lo84+8weKaMuSWirKuWTc
ENL659OxV/OZu0Sqp23ICtkH2sKURVmUeSxtWvTZ913vEdZ19iRKSnB9kz98RX7xTxgESTxzVGlx
u6sjLVnEBUdotr5bkN7kBH9EYXdCT0TiEF9762dChoZ2EWDa9c62u5MAi72kKK49e3HOJ0/YV9ew
i5fDNHBUFVusv2b1RTFEjyTtY9Iv8L1vnq7Pn+qNTSnlw6pNrarDnryJUBaM2Fo4ldMj3UFxN9vJ
tBSaqlGWByi4Zxj6gecVD2jACzVpAU5Q4VL6VJ/qzwGdKWk1M1BAXf7Iejaa2IG0MmM/kcqe7yb0
qr227BNEuxD9CpY3335ZtK6obdu+K3JmBDZcC28gQLXGCK+ro6CKB1gC9L7PONk/0Y2yJ3B6UKc5
rt6REN2NcqFYgit0wWSsHFDnKpx2Y3z2ypPMu4nBw4wz3BgS/tFMwwBQhOSOhyHdVzPwWTmKLbrn
vRnY094KZdBWQGeAwQF+DtHGEzvOOooZ2Ojigd9QAMau2xsgw7K8bc/b6ZgrSpqrvZe4S6r54nDh
AHfzYfqhWcav0pqUnB/BhzyuNeVquQ+W27JebsnBL1WtpKrd3mI8UsRggbyGr85Hcxka/Ojtxlp8
hL3c3UeqK+w9Fi4nXpwubStMUnniYWWo2KvGITyGY0vJkWR68d5rlL8tvOcwazR2MPSNNdwI+JvR
AmQsCByDYm3Ln73MQxTi+49jtY/ABQ0Gu1GHhvpfGSluyYKNnisBiJXiqRvqEEtMFnCR17zSA1pP
ipKBUzRtAZI7TY9u/7H+ib/MvWPiVj/3lixrwAr2LjxoPdH/TrjWhC+QaZ0E6JswdIPo6hC/5gBc
vcbD+oFnqt3RjaD58LuwX4MQeO/oNbjd/PTyr5/ge6Xudju34wYNgD0zJnzBIJkfDF02B5R4z5Zn
2o4ztDrfXC06bAEVLC+WCUl4x16o3yX6DVSOpf/5j0jCMOXmPmE33Ahk7eAzsVW8R13DarVd6qn4
H7j+dJ9Yj1wT0C5+b5z44xnqfAHLmbaYrwk3LPUrfX2yGZ6+oWWbm5J2Q9HAfLlKW44hNeUgoAc5
+CLl8CbjNB5iSjfI0Q1qdgvACbNsZnYeOFTHs1nmKiaV1r2yHNO231APWo4MdG7/K/5rYdap5mmW
3P1VG1UpB3uPjDa4pI5NPU2muRjq16OajWJpl7Q+jLLHZVROzmc16p57WVLlbsoCTiY6foWWReFT
R23XOhtgSkj7tgdCHfZHgij9DYOTqDrRXClv0i5tW4R5yu1QdocnRFY1ZtnQfvHDO0JsMWl+BeRS
JtxmK2MCaWQARm6FqbDU52GEbyBFg//STL0+VhtoxCpOE/P6v5rSz7hEoguugKEUFVnClX3bel4+
SUT4rLhWlp+KklrV1bv/GUV/RjUax/UKorITHsK0Y4HcgDcBL1WTEEG/EEzjwlhNQcxAjlIFneHr
6fb1x7mz75Bn1m+GA0tk4ZHB4P3wlZ35p4oYjggQQh7sQtNC0ndtNgF7VopumMaPlowesHQ8z4l9
jr4EKpxEOyNXQvoqCojngs+Oi3MuxnxNPznUXm/1hPVXfUjL0870NIAM0ey0Jl16dwFW3Bdxar4p
QhkBljb7DjBfTlZ9hDLxdvtsyUx/Af2evOgbhwGN442icLBX0s2qPXmOms7hrKnsvxG/d/yxb+Me
pWAOQz/VPqgZh7wl2tgTMhbgOfmWNezXZPfVCwVWcsixmr3ls5IVlIN5mZrQUydZ4V2XdMK1FkqU
0k7d5kaUKyys9enxCLmM682NT3o+g9HGlWMoX83RCwsyvvpFKEi8uJHZtI78bpfXsutenzXDO/kr
RXGx0r8S6pKfBnN0n9mbr/ggROJWQ77awfZqWKNHjrmNaRPnyDd2/A7hdL1yzxyVthl/zsAMn54Q
ieUU+SP8tGEdiJTVq7QTeSZIy6lCfhfnWZFVlqUzm/zqU/Dwd1GelLkvoHO3WfYN/vWbmzxPqtLd
xxPkk3MMY/9MAw3a/fHCpVHY3Z678hozt8R930OrHShH2Hx+8x4KdFfpIrYg50VXkq+Mo4oQ6rHv
r0ysISF9uYJBjv+cOjb8Tc8x9cenGPpKMYGv1IIkECPSqZI9Qo8B9AyFBT5d/ZruJcsuoHYBhntb
CkGDlmXEBGHWd7AKNLg3d6ChN0iwOMohxd1Gq3qCiPuqUTbnVGyK7ZQqURmDsnBN0O1pdZYjCpjl
Gx74yAFZLlzCWOA6ZlMUsOoESiGR5VszNFbdDVcy6NB1cd6FSyIfWw2Zdes/ZbgU4w/XDGWw0uoi
7NzrnSsF74LdpzobhaCkEGDb/HzNcJl59FzR0ReRQ+SZrzf6MOXENSvYW92Lazlln/omv3M6F5Cn
0kV4rerTXmb8D7zl+Iy/Z5MJ6Tjan+PY2lq2TArQc92EX6grXllmifkzwaIDSbZaStL+tCu/5rbj
Dpi5lad9T3Jpv2UszcersnFouU+BqezV/RGIoZozm9pi396kxqXw0wXaM2Ss+CxddyRjhMCu3r85
QXFicgsVZSnpInK3lTBHW6Y+s7YO/Nc3Ch4F2l4mbbBF3vD7kgC0D9BdMn765NQu9bQNKWEaI5Pf
VRVHH9L4gIlDtykPrZQPMMvPOH2JNCPbsxGy7e9jJAdq6BtEfTYwhAgd3KqPJx5H1VnJqbFo21+g
272xK6DWf2gacMxdUliN/R+l0GVNP0zBvClO+Qai/WMw9iA8ElEIAuWqu+S+Fu40yOVqt9Pb/MG5
H4RZCdkLqjeFfLk//JNUuBwW16WwNQ+s7ig3cGyPEJmF/XytUUXk95MSLnxGPJnMd9SJntXMAv3R
5E+g1BaZFPc3ayyOsnaIEXgkHUoLd7IYz3aGM9guoM4Poe8M3nyacaoXEfv5a/+Dzn4zwFJj/AU+
ah/4K+Yj82qCNb2IvHOPpxXWvm4F+QhlNAA07hS6dn+UBN1adAgu9MdzKPw7a7as4UZhQ/5GhC50
t1+RXasbdfhvMcE8nC+MKrmEbjlfTnyL98a+6XXclynG6+TADmt5GwIL4yX8D+8z84OJwA/eyBPN
g9sirbT8IBuut3I8wVUAU8UMIDHdp3vvhZm+uhTu3UXqxhIgz4cIIuVZG0M8qu7GLR+enn5XytWW
rbBjE5nRqgwTOm/3139pT4TgWNvJFL69URkzi6LHI0Brs79FsQrtz2JYaRD0tijA9UWzxAhAsDS+
/2idwTizwmBEccJdEVUr4wV2DrzSGVPZ4cPjE2ADUJso2ND/2qKxU6PmqgFeXHjwiVSDsS0bhC8D
IHb/G5Xr65G+OFWdDh0jutd5PnCputF8Cf5WJb3O2MxA3fDEU6TKko/dLSMYOi//PKpGb4zunpW8
L24A5/4FCPmDfwpd0mRIYOID3GZynfR1T/mhdcWsChsZie3mFAAWmGiSXitKLsgBk2sopSlc/aSN
R6KF7RmXuzLBTnAZNEbNqLHyhb0n0NkgcOmreSMp3EIlWZY2/p3WxWwHmnKnrfc3WKIsWxwjeMK7
hNun+YnEjARcKCXYi0cGn3ips3ahmbXQeT8WpNN4TT3JIb2OGcDkDIIupMhLNOXM18b9/odqAMFY
+ugxovNQrIt7l+O2bL05iMiBeGiQqYBGH7yskxTK7lbyMVXGeI/vX2zMsKSukys211aC2reSSy+Q
ykcTPWgsTxVCa7G9oTBB+aZ4fOuyDbpOzBEE/N3E5EwXro4aH0nZh8FTKZQfHi0cP9w3/kb6JUYV
vULDTO+t82mf25jB6lcxoEANIwQh26Fl8Tk/3wIaqpi1STYWZhwwz1m5GUPSlALCHwvIr6jSaJ6F
Nkhz0GbeQzBqaahrJJudWzuZhKYGZnSTojx1XABzgd45CZIgamWxf2KirK5TG9HbCppK5o8APnrR
QFfMM1YYUXgTa/VjtTpIrW7DoyvlQOQOLWBKevvhfjkga8ye+Bv0VjhRDW3T00OF0dWTmUN3Cq7N
OX5uIh6rSJwle2Dr+d3MtBVQm0+Ktr2Het2WvaKuVEDKjpVsh9ZR2iPLIGZ+Ax2gfBxybZGeuDp8
Lv0zThtDYshhfn7rc8qsHDPAk0/SkXuwQ8BwPgXw2QloWZA4qJMRFPIECKv+f/yzRfQIsZbQVcwH
DBZlKGDi0nVu78PK1yUWS7z+tK9Plato6Hm2qW+IewFAyoMi7xGD0Ipf3nCuI1GIWNeWihYJMzhK
6GRL7xEH6mKpzewiVPnyCAkjkztglXnfuWYDSJQGyYOlnb2FoHapwr+9V/ViWvLXwYs0IZY8VB6F
BK/hdPxbxOTNRgaDvE0T/UKiqCPfN0WiXnhjEyLDK/jaSjdqIXnTpgymkNXg5C3ugfeikN14dRat
kGtj/l/MkurZ6u9G7XYdZVaVPT7lOsBgHjHU5khe24qKWnRn31Jm9uQJFoAIvoBom5bZwhX5zb1J
hcYq2qxiQLXw3IIAvQ27Ikgu9jk5tM8H0UwfAQl3XE8LiDNqzk2oVZcFhMBtSeaZ43yGXVsLPP4F
foieHWFxbo2ZvW8ISZTzFrDzZQdR3gQ0KXC4hWqp2oJd7gBGXFe44lq8RXcl2UrWTYhzgh8hCfrt
bCZzABzVlWSZLH9yRWYhKI5IjQuObFZg9q+cpo8UXwpvxO3K+zgVWlo2M6mq25C9vwgBf3vPXeaX
D/zhfo8dkJ4eX2g5dWLC03mRekKTAhBvLV1CQHyr1vxdVlufC6po88n5xtNTu4PAhx7fKUZhsH7C
iyi1P/jVI3rXZIMuu0gQoAaiPHlmKxxL8K+lDQMVXokhH5S4qzKP5NAQrDUZr5uyveDF5ilV+ijq
wQ05O2iWoj5iISoIwGunva3r8xsSfLTAb4o3gA8JWMIThPmanO2t4XxoP25b8uujsyV3uOD/xmnE
axRN7C7UqC+4GqO34KzWJ31z7eA7i/qGLGx9zdq7k9/E/TDMexq0JaYBntZ1X6VGoHwLUHjJn5s2
qgEATbJFJqUB8wvaUH/pBoV9AtjK/9ayw9+1AtVWnZjklKuEbYZ2JgNgld4yuzqHvO+nvGOIVuK1
xv0gQq5ucFBxEZ8OCNjN8ybULfkp5IaCkWUjUGozr5/YMsisbEKv8dhcTrLV+tN1rZik5y0tKPLM
QjfFvOUYjjX31BAFBPMIxIcHhCJ7lXTvyYABqhqzBGDM5xr8ZOjEXo5i0NXMzDTavTmdXUOA0M/T
LjY/2uc+i76tp5hUdHSbnvoWz6cmSkOhrS5DA5yNc2Z8+qu4oaYoQ630CX7So/qjQxUzkoSQ1Cmu
U78LChZGeD9s54w/PTDzaSJvXPWenrpEb5+75fGp50SsRtsLreUj9tJyyIqEQi+oFsf1/x7zBsIp
ELJmMUgNESiCssAFr3G8KtizlgFs5plJCMsTPa5hRrYbmh0H5uHevQzej693VvSvqzvGSiWkNQ91
27T6gDdYkp/lbou+tMXGXYcn+6Ec3/wHez8M4+SDsbbK47nK4FTB4AmKiqVeT6FhhE7Q7A4c0VUf
JnjogKgMyF62iidoqCeevun6u2F9lyUgExjPllGUM7JWI77JkUQL8cFMguTOseay29Byp/9XIje3
Hl7C9EBQPMkbHynqjyeiRA50CI6UDBCaGZzEr3UquOOrK4pOdGpCjtWJNELzVs+UnoM02NdexuEa
bg6/jVsWKAuKZhMWn8Uh/r0wJqhXHAa9MPHjOynMVxJp5oyerNZb5A4NelWP+keP0lriQ3NBlPYv
7mkFTNczJMxSofCOZZs2SmI7nlAzhi6jN/+yc4SrYGSj7byDMLAgBT27blrnWkK+SP+h4rkGrEfx
YhIlTdfbhDpzh52KLhurc6EcV6mnd3SgN+rEzpOJNEvrB4y8bihwu8xD92/ypxM30CpwqNtY1g7l
28p1EAZfM6iFrHKY2xbH+ise/1IXdbsfhLKVH/znCBmt5ovd2vvrrpmLOdDwh1jNIq7t3eQ06jFL
ccrG5MNFltcCX0zp8S98GASO0h/rPcWKRMve7dtm51EzMV6ghEbJKClnEzDdSAqBwdW9+2kyc0I5
YN/hE0QV11OmFfUlThYO8otixOUaygHuMVcIIcVGvEjhN4ujzIGgvp8II/z6VXKE/M74SJkFigtQ
69aT6yxvxw5aLkAASR+v5YHDOh3ocr2HRX6oWIgG2lJSJEzydzAbjJ1Hdx0shVOS3ki96HKAWBUE
syko5wmizC8D0IO/SqgIVctVvOQ9rcHXOq4rnHGLEyjNhtUjg/9n8grRX6CI99jo2JirCUWMKPex
ZSVKYsw6pGux8AkqCxncvisgjXGJGSNXGL8+EJ0xNeTJjcVFt7jthbPoeGmwVI9HGhvuSPC+CdgD
dpGvRmSXebiC35nVShSBJ9sB3UlQewYT/5NTIr/hBvKB5Es5L7SajmOiHdsWHQGfKRLW3unXxeRz
WQumkT3Sg7zSKFQGVCQ23SwvsK7Enj8D4T2RU4wWuqpTUjwfxsrao04cUYl9XSC5IzAIsh5Skv5G
dOP4hYZA3YIG/pb1zunv1Vy/qkzqQsXpz/ksIuemFpd7NeueqzRjQQygqAv6WFugsB+7Fn9BJelL
QDXjmeFDYb32HH40A1g4801mgLTzKU/31nP6WMw2PzZEInfakN6HSXjp36TATAZm8s8ojpkRowQv
nk2pBVimxahRS88JKu1muaOhhtEHa6OTibrJZqrM0Ad3XVIyeD3iOBALVV+UYmXMurbSQ0BiqIB6
Lrw7IYDZJ/xFf8+DYYxYXMNznXW9kAiir3x31QKSamQ7RYGmqQMWmzp6zKYinlPNRnF3/vkHpHHB
dp5gz8rr08GrbA9jlL1vd75COh4TGBTn1XakS+CPJB7Dxof7kuJ0obWEaWtt1ALzGJf0P2BK/r/x
5fTcNbOxPfb0gzWp89NYe0CyK+QRONhsaC0kTch99vfERjO2zsIE0omPNU8RKVp+VxcScJMo7PGu
HZy1ZHxNsBToj2BiY6pIQENR410OjttTHIfud6U7v68l5PhQ0FZ9GtnH1Ja1r+SeSpAzd2lFRii9
4EqDaPJXqzOHeXLIfgB0779uVZemf3tuayojE4vMLzKAuk0gnmcl0jXz/FDAgOCX1iwlTy7oHMhs
JG6deRbogvEKv72Wd0L3Tg04H5jsi+wZCFAeAP6RNVi1Eba2QiubhnLE882rd7+z3fFBHF5/3z43
7s9Zna7zV6xfR3Q20xZY7Pi5crk45kAXfLZneeRY7x4xjIWGajFBK5buCDJr4KDLrozdM2WOz95B
w4jxZQmZFaTj+DiUIHgUyY8refEw5Fcmo3cf2NAv057LrLIDvxC6u6NeWANVQpqt+eorFsrKAhQH
laWGxkdk0+s6mLpYWxDAm6Goy2uvcxeU1Lqb7QyBKyILZ2PeC1HnRFKAS2+hvDV6XUBBwmWIUZlS
dRgIdWGB5eKargERum/97waX0rC5dc+tGGgWGLfyVCHjAlyLNzszrQzV1cRIxbzRaB0CYkOf+sPu
l2xEimRWF4S2DIfF7o4xlpMhnOKwXNIJFFpTOG1gWp527YjY/mHmO6ux2WTVKvrNabTFNIZUckS+
sI323EKBcyZLIowVwObw+hSm6LqSszHNf/hoAiE2zvtALz38yelvXE6lFt8sXRzVit9eUYDEztZF
cUbonKxb9flpHbh/Y9yl9F3q4Bp9LyhO+XLc/cL8/CjTngaQ4TXuaizYHbpOEIistI7HTi78/usR
MSQSrljqktf3G0/UTh7+sXXEFOGTXAxZ+rJC2CTaGYNL8Yb29bvdxdSIRmoZHNtrN3mdB0XG2Vak
aYFnVhw3NLfxMZPHIF+s8uhZA+iq08S0V+yTVZElN0NtB7DhmnDgjm0pKDmC+L+ddgRDEsYsmkg1
YMiGSsFn6AeOUPNpdzRf/IWb+7hiVptMXFpLBcDm2wSg7iBGc9Jn5oPzCzkgk7bd/fJwVzH98k8f
luuLbEzYMhHudnMd4dW77fyfGjRWg03h4zI0LiAAJbsCehemkCUy/YwaRwttGvE8i4Dwn8I+VCwg
rCyZ1b6j3OSCMUvNRD5cKt3QIInWz2O1PMNhp91AOyqMhdoEGpuAo3sf/6o3JTRxVkxfZKwHYB1I
Ej/ifdoLZpyjt4/jKmOVWTucM9gcQ76euQJCMT7bAEm+Khe6ctsuy7xjjT3mCDu07FSVkaqjjAw+
95RcK+6oOdn9QBbDR2cqiNAaFPmR1SoHhMmGw7Qz/qJKijWsOSs3M1EU/cipMCtrTFfrE98NiGbY
z04G8CYnkAA9ebxMm14G9hZf/tPpG1CScy+dCN7pHNa9XPY/Zqz3seuaQ7Z/k1RUROXe+uW+MDTo
2uAqSu7EUT3oGtDg3pMRqyAQWvLCddYr8/q5Qw9ftwdO8fF4tkRfSZwzyU/Uu+fOK9mH3gwvLQol
UhF3iTB6DHjqI7CMCoIKJi4l7FIKUifWWrPbh+wCsdmnW0BGvS4XpbOaw/6Ao5Jkb1FxlgbHEO1j
uG7Z3HJCCnV22QDfDUrbH2QnDkkfUQsFLQI3/xwWSqgOCe1RUoSclU38sdXEkcrjLJK6alRQ7nTx
5yIR48QGw5yUmNIjH5sV83yapZkSPvxJeAlbFTYI3lZgQi9/kjmT6h5gkvC93u8gTGtwWw7LUtTd
vy2HYTvEjeuO6XacrDMG6fD+jO+/2aDQOeIdgSJE4cwJHQzmI2XLPnGPesQHS6ksFyPXoq4xuleM
ZAgtQFM2r6OR5RE3mdn8F53XBgnj9Fv4dykLVG9Q2tLypo28NKvtbihYiIl7cB7sUta44h03CSv8
zGn7G0HCJfCkkq1hps9R6haykO2JlvzA2cAuAbmQbJxsHtFBUBcKLicHU+nRkd5J8ZKh12JjY1nD
gBuqm6slXmpXpoSuzXOO+B4qwTPJg7sUulIqnn5OYroHD+gQU00bzVfA7/CnSTQ9EpQGSDfHJZZb
FrH5svoVZnMBdPc1T2Yx94PhxkVVJptseqA60a0tqXlbDzUScEIfm7ywvKNF0jB+Ejts4YUtYDN4
9WFoxH0bljEXEs1I8MlMeDRZ1xHirSgmpod8ur6x4GwLoumj2LDCVS8jAgsLRRXJ3Uqq+D716l9X
9Ab/tVbMFVjNY2RxwmbzRa0+atRs4iq2KMJuLqIbYBhIGlMWONBwMgmPjaDVz/LUKcgNPR/WW3Rg
iFSibFVznDJpXkgqERsmbWxBGnuEt3J0VpgbsGi9A0pNaVEEPXO7FvMDTox23lDZ63/xwt3fKYf7
YSz9Wk1ErTWg3kaFNWx9X45IBybJRIa/c1OATSS1Nn8GOFM6g9m1wtBcJ46IDHfZdXvFv1OCEF93
s95c2ayonvWoe8zqs6OUNJskEXnVgPFU/TKRZBeabpSCA+4jx8F1j+H0yQURUqSjQGyrk5h/Ct/2
jrZyulI28LE8edSr4ycApi7OrSKmyPx9Q28cxwU6lxaqmtH82pjySPt9HnynJqjNTLiEDi+FNLUt
GosKrI30Lf8qiBI8TT1MHERjN4ZLgCsNQRw/oHrmzBMxXaUFtVOCJbqc8npRf/SXrLb3WXynEVTs
tYCEW9SkJ83bJpDdAH1IGMUXFzt131hToryiGvN28JbOcL8qj2iyfMlhj05aonEFMLupDcWIjvBz
JFsKLliOtwABp2jZhmkYcRuRc5I0wRoMPWX6OhHHgen1lWcd66dzJN6fG+L968qc0KkN5Upl6q9q
xZYKJTDi/5C2oQ6Nr+2oFNmTHCUktFpe/yyQZWUW24ybCB668Nb8B+7J3Lsc/zTkUEgjvrv5A1Nd
vHNHik3/cyW+2jluW8YTc7w5Mj971CCp1FwlUgDDpW9nVU18xaoPRSVMZMH/sWmLCpuGbyiDbonB
337GRmjHnXaxEbyAWTMZC4A4rk1N92Z2VL3Riujc1J0xBAwJrSaRuO3hm1zePnyFVCKrr8Ql5HcB
xDIJiFrpmj6sseyL4FLj5/jnNwDMGAaeZIoRiQOe8+HOuUMTGtick+MuHBM6VA11H9GHkv0XliiQ
ltaB38zrmy/2Jmtq296PzfLYbceqOGpsjjhLBn44SiH91jIulohx67nWPwLAVd1IBVqDvB+4GRNF
VBC9kEc6PzRcKw3+yR3eCYFrqxE0Qme3iu95mBcLX4eLNl+YRgtCjEc+oWugfzUAmBgZBjgciiFt
xDIHfdQveczllAHeQ37eCyyo6PKo/vAZ6Ltu7HWYZzQqK6skGnuYziMXDAf+GysmbIjLHei4OjV1
wLF4GmWO+uA2JwNtvTxpO8y0JWS6Rt3WHfu5RenBFMiv4F7Bf5dDHWXgqB2fPS/2s0ZZH/y6xByc
5Wf5gU0lMH1YD2dMqe8fqzeDVOzKGgfI9TWZAyJuCeezEozDJHx/m8SIak6C7MI8KJaCVNBch3pw
hqxCg2DG6rZC/E9yCrY9+HnOJ8yyBtndwPREFT4Y0T6DGbr517U0KYnzpYIdPKXapx3irm5ZaNI0
rMGUOnelZmSuIUyyihUddxgC/iQpL70bS/XIptZ9xlKnZ8rFCHnq8TbaxL101LCGXqAOrJT5VaMU
KfKsiad+xMP+A13Z50B87vUmzGXWe7sOITCU59gbYim+cnUwmCsjEf3UyIvnHHyWdLavhQWfQRRn
L8BNy3srEnHUCWfLar8+tMWB3XHGJvSG2GrIi1otIEAyIca1J1eZFOX33Jy+k9arhMnDwxOXau0y
urQ6Pyajk614RnYy7JKEmW3Zd6TN1Voh9J9nG3Eo9lxO1OQFaDbzHBeuLqs4mL72rO/w/DO4IAtv
JPMdH5iMtSWy9eIDLLvMO08U2SMzRrqZ9nMjTxlnipf/RKfW601Pdo/ZeIrEmcmixCCX40+Hny5c
Xu3haC8pm1qAnBBbL9pVRi9nJKB2MrEVtjRlG8sUQJc9CS36Npr18gQNqGhYeLgZVKlmQf7J9WR2
+qdWwyK7HOKxB4lxYGnCpHfOaHhl4Wssh5v/zVeBTOjGO2wjTEWj3ZCfW2KXBUhuTbCMJs9P77vb
i6wkAAlnUIAMSGJeaqkSjbCUlGaWE5M91joaSoNmWYVbqJnblwevFdoRQt252uLb6je5QiB3F1pJ
m5FrV6+cEeUV4TbeA9KIoYxmDuOMgtHDaL79OFpuVPR6YqHLS4eVwHiKyHFzdebMZ2/s4IMzQXg1
mCMySjHWBP2eYQejtwdNeSTexKDq1Z03hMMRZZY5lKglCbCOH5GS36Ipx7Q+qF+ri41AUuyc+JKh
AEoYNjf3YnaJ/k6DKNGLKF/wuD0pG5g5LT2TQ8h/gCHo9fWYkVfhMLzfpmVvfYnMR7f3cNnrx4uV
ZzCog5cqhVxfc9xogjksmCnUv4QM4bWuTFN4hMsGKoXD5gu49y6BsYFfwRjs+kjZOedLY+LfAbml
HLm4nPe5m9vBH9f3k/Eb2cwLv9+efnRfjKJxO5wP1S5tdr1mwTOeGoPcZl5J+7dM2Q6Ef05y1u+w
RQvqMwPG0fjzAOWYBZODxpTNrausYUPIy7pXBRFZ4ZsQkLXt/9dZ0PfD1SGBhMugZlaimcjDbajh
NByPDR3g8CiFVde3+mDiTIHIUKDZ9m5CXiXNGTsr3nDPSbm2lvZUF0EVqX6IDvKkKS31mqR2wgSk
ysL0kgrhEgahu1jjNn4essGJQjLAAIAYuCZPqlACOW2s01yHNoDKT8LozNoLTHvoeiS6suMLPcnE
ybyIpRMZZX5p+YV6uxNBUeycC6tJk3Uz185eCpO219jqw0lwKO4h7V8taBQao2UJ9f0a+vlr9Epc
XRpMr9lvRC2OlaGVhTtqyfsOyaWLUfnF45UppF805XTzfhepCcSEZnb9XtQj/anO+93XZJB4VpMU
3mh1/zJa9E+PlUboiulBsFFrK7ZIhjTIuU6B76Y0cDS9QjKNWmiEdTz7rE2iMNOvjV+BjmtBC9qd
JAquWXAz85NRTAIbL7Nnv/KLavW8zMZ7grAjuzuP3JkrCkebXKN3zBnNgCqwP+jrFQHu1Ghjd1UM
rgDngPHUWs3+/VCi1O+WiCgqSnyN+MrsjRxj48ptys6GvSAMqWLkH+69GgV2Oabsdf6ZHLJbm/81
PrmEuH8EBCPEitE1DVLsgGoEhftuz2fhQth+qzl3GRzVTy+QoNwIm/RcrTyHG+WIYVUF7OHorlNs
f/woWh6aGlpXwv4/yseF6/U6EchLYTzFcA62u6hBwE3dKel5hwoe6rKgjncfG8kzx0ELlj/IwdWb
IzBtinVf5DAU17kvkzWtoOyPr8fu18/EQBPw+YfU2AZeMZKstaRUrFKx5DasNIcLcOS9d6vHnEX2
DaNTCD4M/xZI9Bc9HpQUbdiARuVY5slIQvzRnXCZYXuuyb5kZ9CxlLEKCyi4oXo2P/dnV7hLb0cf
O6SF3LnnT0nevV/CYSB8xh7YkK/rWc++P7L44gJ8/Uq33boK0UrAakfs+t6BkSCpRBmb8xaFQvMU
jry7JVp5lBKPCZUG5DJdoWoesjYFmfsOwzcvUxVDzLtfVuKVAHS7pvn6LsMZ3UZFPc3Enn+4X8wR
1fn252SRLW7+E+LCvWKJ96Fp85Sod3zTK0uH6p6Rf4ks9ToUxYaGXEiKFDf7781FtIpm69Xn0YUb
43faaF5vZYZD81RHddEuR6FQeaLhhYK+t0r/LVvJfhtd3CBfke1YQdqbH8+WTDIX3+sUueu6EYJV
4y/of+8fc0mrmKctJOC6RyeqaFIpCApeNQQ666LlrO8D6GRtQEY6BegKihIHUZ6wmv5vZ+cEsk2C
f4Yjn93cImf7Q6zmaWk/10Sto9bNu6sF9/U3qkyE5lpf/bKiKX6G/rTkD3SmqISQ3HAGH9YUqx9F
u0Txz/f4RqIpZugi/Sdeo8gudJCSEhL+hp2dP8hEEmUGxzz8ysP25Xm4gqnAB8L//AtHIQXkf8o3
xEmHpw+G6SaqNSYKRRWhbMKjbvUzqx9zlS+VKaR0YPODHzCccqY1Z7D6E+LVkfXOQymwv5ND8WxH
q+FcIJcSTL9jN4DpLvWmySJQefakaS21AHGjsFCIl36Hlv5YiskcA3ttk1XiR9PGAAzXXOyrrnBj
ZJDapUhjGNcOpMa3EaoXcs05Dg8aFDEdXtsyLmTM1P66Ts24DKLDkVlDMCs1j34ndf39ZbmUulA1
MwSgIoZyLj2soAlIeIlE2Cqq+qbiXfeZafSrGILckI+E3gTNsWJvii7B/BZX9HSAbB2NPw56d7t/
bq3R+1bAI/zwqIdHw1sQfeVYWQp1nIi6MEZ2U50L7aEDDf6uNRAv5MaUIafeyK5rx4mtT6lkddXg
OHoHSR+2lL/NqL6QuFfxotoYKqN4K2ups/tlwpXC0B06OwALDaZYWK+pEAXWt9HK9jHeLpgT+WLB
pE7HEnPFrvzmTbVHY1y5I5OX0FqmfOfp8NbLcCiJkiLWXIAEkoxYu5UzTYgmcNtHiJGnizHl1nv8
b6/Cif9rvpK8TI+wr8oFtj4rtThzAi99zXbr9XzCnt+c1CR9dmtjegckD4Hpviqim3bFTYyJY2D2
1PTwDgKcJoiANBA5lBHCg+KQEvksF70ix5Kj2PhxCmRcyfmlyLAKV30fbMOlWvEjDj3IHVrpDgsu
fVzHdw/lTR4sm5OEnE8dD6fAoYKG/eJYltJLBN+6Zv0KpSTGef6zvlpPELyeXrSSXYOUYv7euEb7
ZxcztqX4XoRv4Lftpx644cOO8K8DL9dkuwrsL4I8HnBZPC7ZYNxAgmbpvxJdji/ypykG9rse6hib
w7swhRyMeDOSa/VRJFQJGGthGOYOaNRpxxdouUBTRckMhs1NLvBErDpPkeDFZEiF4s4GTH43Xce3
tE82KVfuhAcJ8Hj2DrUCfBxPrUqje350+QghOKQKOdbrIBw5UiZ3/i4iNkNDo3gX/uIxVdKMaDrS
v7sD2lFredw1ZA3PtGwBCmC6FUuzYwvVpTMzc9qGlj7ZXDs66+0aFM5J5icQEqV0xBYtg6nMxRvx
zDlKGU3hYd4ce85Kw/yZdfXjtV5iSOPB50PlHGvgp6qfLQAjDdLHMiWLiJmT64IPLPg831uZmwZs
BtL4bHzQ8IvuS974EFvmouZ85qRNWhTGk1LOnOKRI0tEw/3FGIXBND4tnD8uSrc1IeQwv1NnpZDk
Bim8SfsWPSO2AFWSzPKFgBykUUdcAQIAbmScOE3Xv5cZwAHMGUCy1ov+f2dJYDO1FzBaIG8BcKPa
2T/L8BH6JShB/XBpSdwh2nN3kwhEWbGHe8eRapVLEAT0OvReEJntHF8FaTj4x/Ahz/bS0NvviX+s
fBGgX89jmkCWBdrTK8ggek0/oPbA8uGsgFk1b9iulIvmMDhRu08u7ajz8wrIquwpbQu98UeWvEic
KO3Kzh8m2Xq9IiMdPlHA60QlTfgd9niP5GMkjWTNaZj+HtfdY9B91CmUYi3Zz24TLggLxnpFu4mK
S6cdC8k/2d7xd2b+79YC+7ruG4TcaolZdP/tRNq8t66VRD2pBVoE+/s41Ah22OVEbiyv+VUTB+ac
60PhWbxlAckCYz6zxemalQ3wJeYmJ5b7h72EFQ0VyAIiSKdmcRZ5nOa83lXrcLr/vVgN+evF7N3x
BErc6pe7e6E5Ecic0iFE533YL6EeCC7jXb3pXFBNwMZU74qGiHIT58iQjTrKgipMSrtUYbfV9IID
/HLGSUmfm3MebWTRltiXyREi7a43CtHw98JnfRPrJ8BYOd7KZeEhbdKfAywCp+OkbiwP6pvlgZmw
/PfVdMWNHLHL/15wK4E+qcXCjtII8O+FoQAE3zpGzF9b8aBQKQoSoSZI5XibaXym35yLQ6jNCKtL
uDdtct/o75PkH0pB5hUKt90k6j3G7C08HP01zBYIts8ev0Ya1T0+zHqKx6VrvgjH9IkVABvmJhr+
CxC7VCozZR+PxqXrGygVnMDlGU4UCZckxh4A/CmuRHLh2fWGt+C3KYn2l+n7KuJT6iH+DyP+iCh6
+zXfQD6fyfrt9RwEOUURYEIh5N3cQQY5eTC9ZqDu+cWGd67k8VpfbuTNgPbslVxy1m45o3Ml/b0P
/16rpPOA9jHWHPjUJ+QhlE7OrczMbbKr8hZgA2sNhDQzimPHxjOas2ZVbQFuBzVfOqZlBwdgidAw
0B8750xEfWWNVqxB7BWnyvg7/qQpF/ifeBmLyKOIJmdCp2esHd4inYfAxK9GfW2rzq88tZoPJMw9
wmJc/3mMLZN/NBi5I7/NcpUKTqLrtV7hBnwbJJH5YXmeFRvc9PQjm1Hntu++aXpNUx4GaiVc9pSQ
Elphv35OTyNWUEsMuW9q9y2SLLegyzKrZdQIchZKML2Pxnli6rEha7sfrO7eOcuuAiSkNLUsS0Bz
gJalb64mLbQH9Y8OtZTwFk8O6iZp4tE77E9T1uFBypjcuYw4BKvyDvF10II+oXvi93YUcfXxydA9
TTz/bcGy82nwIt2Itbb2wnYggkvpi11lp+4IdsoZVyIrLEuaxET5/PNo9In4FctHc3ImhVJwjrBQ
+MbDxZXN84OoXNsgGcIh2fMmT0/q6rJAZUt/RKSe1peYAIaFckW1PdvID7kYfs2KPa+Qa2waESOJ
yzqQwRpd1bqdf125mZQQ4AS/RKwghrTYZ6kEOqqv03qJFwlonAfAsmkXjjmDhqSx99RJmXbUCTIC
xcwMGsbLiI7HEwVCd8LYYRmqGnjKrMAnih/N0AV0C2E2CQLNWiRM9vnAXNwVy/YNHEZJoaObMm9m
c1HUbGr3K+OgVMVp3IoqZFT2I2C2f4sPwD1905vwef0xqHDEJIiWTHzzjQjNrkicfINnIiQi7ArU
gq8bOWUgEPX4WJj0O9BzoWq92yvvxW6BUXR0Cya12C40xcrU/G+r5LhskBvO1oINYm2TcLiju0kI
HxsjVRrvbrzFGkUy3i7NEodsznBUqS3OL9bTXzR/QAW0w5yk72XB372UCWI5gQ2NAwX/X9rqEbWo
y+DbyUeahqcV+zeo6hMgjIoVCqi8aH9D9Ls1/c0S5kWItPChibDu9UaJwymrtaRUkcBH1A2wvOi2
N/or91J/zKDW7M+/cVC4rbxAMDdPEBCwBHy+Xgb8x6YFFa6u8QOYv1dYQIQu316yhM+Oq8jzZFAc
BhIopStFkuVmYX5xroHChEyUa5YHPD+7OTJvORN31L0vQq8Ex4Lh9bk6c4KWpYx7lCXpWk6vSEtP
bTJFQ972Bj9OAxSg067q/mNwH35HWIEJriKRNUP0hMggV7E0lpMwLOaRUHBR4FoEyum/FM2NqHz7
XMXPKDW7z7Q7ccmGIIRtxeP4j7Hwd8F8swy/M3dGRthhBSj6W4PWnXjGL+JGiieJi1qGPVCbYSSJ
xCvuTWhsm9K8jyaYhH8dwSTGDw2vWRVAsquOUkHVGXn4RN674asHKOomhhN03NyPnNYZEbwCaqPF
RKNfKgiTgycrOH80yHQflZRwOXLYRLplFq2wEYQ+zYB8Xc4nCUs/YEuRe90MHxPT0tosHWYeS/BS
FtJXiE0T1VI4Sv3CiIzrsx6h19iwawuRK2NEo8cEZoW3jM0/EkvaXubgV+sTXGiO0MacW1d3ivOz
8wiK8fKF/Xwk5y9R4rbeOraUv+8teOsjypnW0zVL7+FascHexmZGuq+npZEpI6GuhJWrx399E6vh
C35t4fR3uSKSwDIpmwShGKUWxmiQ9LlVnqNoiXswsxC/tqTmu+VZBxcPvOjejRZZtxRMgqupFIwM
gCD0gWeqSxkahScuTgUVBryBw98xe10GXhjmoxWd2wiZ4hgRqmURgtZ8Vh6Alu88NhwL/YOl9MoB
nF79iWGNku+VDP/KxnITVKCHn28xre1A+dkZoTm0OBt4dMLgNLzWJTRZPNOnWh3pz+G0VuoMDWUV
1c0drIpUOT+71UmqekZJ7DFjyksBgdARFuFY4+hfMV0aGHyYUV9W3eG4PPB7iZXbR3qP/hQF6uiR
dz2XzbEQHSPwEiY6yGdV2izTslz4Pyp+ExCmklZGuGSL8PvUAmBqwV9OVZlQBnDFyMyuzZiXEfjE
iGrYDwAUBRNCU3K9AFo4yHqCZFvza0I+RdVjnCBpiNJTFVX2qV9Q97EryJTN9qORNCsUP5C+QD+8
Xiko+6Vgyg5yEjgZKbF5Bklc+fz5bRrpfjbx0zWK37YdtHTJjC8yAt1/ygjw3PCiKWS239gkHrEI
yp8fPjbxbBVTQcI2GbDGzBNSXIRjq+z0/r+GSzDbUZe17ReAZyWMrU55fI99bOMldR1VsrdCmx6f
lYP3Zuf2iABqe7IhG4LoValNf1AXx3wZDZyAXdQGlGS4lt2wDLrX/zoktr9G5fyFk0Vj0n+r5Fta
p2bKBvVmzF4BTZGPXpIjVwa0/vD347a1fSTAxQppicdINVwzKZnyfYtkYMMtXmg4TnoPL+nMW1gO
2ZgQXvgQ9P2P9l/6gopBPa2xUWSVNDitSI8401v/HPvi8RB7jjmPbHiDtnrNIR4h7WRVDpKaqwHk
eFC8EduO3Aphfp7DVLHYq3610gXVQZH/DnG/a+sBEsUCNyZ8XDNmVLnF7GcDMQxsjKH6ZIL61A4p
kTjg/nvSsdnEFgqDF/4Z6S4EgNJkfT79gXpfjMU/BJv5yyUJ5WTNnqo+LWLH0/SxlyVm/0Uu5TjT
92pqr+mL5GssRcfAyakoEpo6nRaT3FG9DecB8TRnQ8IKkMbeNQ5SFJ0GUxkuUClStQYH0seOmNg2
nqtlyP74jSrzM2YoA1b3GKKmXwyrowcE3ohHF0jBiiRbCU2dyIeXRCqxLmsPZO3Ud4WqZXcMbRFC
oCf8RAORlPnW10bNZkZN6y23reVbldFj1DDEyJ6wH9WGRX/VXYWEU5WaFJlvXMoSCywllaM9ywU1
TRf6nSC+a5TjiluLV2D+l941XKNf+CwVlOCb6KXvKLXZygZBDkkH+8Or9zXf3g2GzFlOrsQCN+f6
qdPCfNo5cj2SgYDQZb3/s7/gSZZq/Un7v5nzgLDbj4tUdBilEqiDEBu2L2VpVa3opmauFpUqVaSe
ovpxeKKH9HjQdzodMZR3xAOLY2JrPgoa8Pkdn+6WSly/X+NRtMrLY2cWl/E2bqzopMiRkWI1Gz3r
9nm85B3bXWddXIselaz5pBDXXul43rQZC3kDmAvCi1R0dPYNSolTSeefI2ce2C8U87KZikLSq0eU
oV0geRsCKdLyZ5/4f8YKequPARb7/iKk7TCJGmazBu1BSU57FjL39t6WLyTqAp5ohA5jDwu4t0Wi
3NBZbZwFycD0o4uPQYH/i6ae+pqw31fqZcJOo6rwEwuV/4XFRNp3+Y4SxS1tq+WHg08QQQqsbAIV
YJWrEZjzf+8VO/xowqm7uori/IhMQi8DeAU5s9UE+9zHttipsQENIdFMt9bYKJ+5UqJ8JINmAKJ6
gYYpeTLgg6EiG9MPykd61sX/+4c88RcLYyEcJjFnRcI9aaLkonY/qc/lbij0ypDXdajswQ1vvylv
fhE0ZeN6BXOyB7m3XV7FI3EoYyl4wrq7alKKYv47KmM57IMCaOUangeeM8wPZZnxeIon5dT06fUz
Sg+92HtKsL9JGkYd5JTPj2oxAZvZqkGtu5JNl7DpvbmMnkkF5CUFYqCtakFAOcleL7XG/vrBPVgs
9lkV/4+KS0AuJUL/2LmrXO9pjlQqAYA3QqKmH6b3jIzIBlNwuzohBjFo81A7+o5cKCD6rii9W3N2
2Fa64lXSWDfcdvdWcaUoCYfkIWF/O6NeRRVuNLCynn/Lb8YVp0v701scUo2mQRP7q5KZq77kU+Qh
yQZrAzGBEOXn/yEYFlUhDw9gMQ7CXboTEhGqeaF566Vu9+oREbWaxlDATwob3X91vL4be+bsw4KB
08SWjnBPtOzprgnDYvwdEN+ThSMB5Df0VeL6CBQDPrpJeZoOAJ1hsosv0FOx7E2CEcR+gRs1U0oz
paBMkgyVgjuKHEVUUjC2A6YRoEUTd3QIn5FgsFePGcWnZ3ro9x7Bbe9Gva9/RZ/onA4Zt/jb6+PX
BpZYyIwRS2jQm7S+IVoyZJVhYfiFlCcQeKCJL4bMR+ClVIZjqnRZ7+GaBORUlgKbRq2XEEzpW613
HpFdPT21GHy/Lpv1joGhWd5v1WUk//dmhu54GBleIZH35rooBl5Ibda2ciTGIgaL9lsG2f7ehoui
f9JBSfBy4+IFTfpyXX5qh6aXZZLESnObPwNBxXV5InGJ2V/oIe+zL4cd26GLm/ya1HK6EGItGXCl
f1g+RGAaKifgJI7CVu1Pg9B6BlO9XpJKRjqxcVpamEFyvJzJHzNAOv9lHrZ/Pp+xvIddhz3Y+XID
H61/l4Db1uhpWmusUip+rQRgdwt1l/dQYsGoG8pYTIVZeS1mLsZttlAo4h1k4A330od6NCcKkXh9
GBctfoEzw/R5yAJSln+FDyAFDoGw9F7pkQSWdimb8ZJiN/A98mzUlhsSVk5G5fgEFbUcDQ7Pojdg
GqdxRg35P6KIlgJbo/Z/GSCCcKrZw4CCFipbIRRqGqpu4+yrZ7bZ+aIyCiot5B5mUEjzQDflmKh1
ga0cLtQptfk2F2FdkWB48WfWfiLLo97HDE+QicwMxIVJzecRgkMT6dh868gOUox/rXUm9F1fJa8P
eH6bbwEu+M9lb/kAWRtrosRHmR4dmMQF8KdMa3w1A8N48c7hlDOjNzXrp0DfajVPjY5WyjSWU3/J
xo5hD9d0/Z3JJiYPBYzG8udWuRXl5fO04N3BmC0x12/dNIMb+EtqyXzPbvpLGDWcHSMHwYciKa1K
+wFkgu01aQ/keF5P1hccZCloddU8I2QN/HXDRzt7OfLp9a+aX4vmHdJX56x6JgJwij86g2y8hOsy
a2ax5GcMI5l70x0+QjJZ/6qm9FSEIGVBAzJz8pJ6qoa117kt7fKkeHqtH6+dc9Y2BT6BbBt37WzQ
dh+jPe2dlS70ET9YiQ4B1+YrzJM3m0Lxam5g0egbRhK/FbpWqW0Q0Xk0DwlrRRoaFLiySQKwF2en
Srfe9DbfHZ21Usv9UZoiUKkJt2SYAGBdhdXzOCR5zVGJKhMevF7c3FrfQUpfLDmgUeiMBco85zoT
204Hyr3QbDSllAwGAuauN+XJS03s5HgRi2HR1hXVRY1bVxYWOrABZpuLvQPuKW3phDoaxFrzT6F+
pFH8COBZa2qG1AECIrCi8zo/ZYs3zg1ubje8XxfLqp3XyNHHvTyA2yYTJNyulB4WzOFcgF8kkAe8
DKQoLXml07MwspDFI+5rk4Z43QLXBYvA5pGFSaX+tJf6Uepqrlz/BVqr6O2wKzrYwWyg70NxnSDi
VJFB70pt2+0BGl3DtDmWcaKli8fUWHbJG5YlailOCzPP857HdwtthQU5jL/ziq6CTnTeDl+rpRMO
FtbWIJCpJO6jGaDS1Wfl4hNxY8XGeMxrNVteHQDUdEclcC1Ot2SNxo+5hd9dvxihTHcUP3PSO15X
gWYI3AE2x/ANWyMJAYSDQR8nLxvSPci5M/+fRVtJCyk6aiYX0t0mdEwCsXJKZ+CXeR9myGnMQBvP
nO0vCqmDjv0+iDSEoDgR6EkXu8xtPISynx3WRiEDWhV4o6C/vAygkll/uMZWIpNy3+MDHwM+fyL0
f8XOua03c1dVGDc2+oTaq1AG+6BrNLo0l8RS90HAbw1axcsjE1yXGsS3XA8eLyTo4SynaB5ev8Cq
TuLAWk3SYwOYVn+GwVuEMI+NFP4AxsDgUEdnMbv5xQilt55E/7Zg8pcUpCQBgS3FazCFyCiFagi2
x6WCb9dmKHpaJba55lAQl68qi9lodjr0rYgzLH+BFlWpXjradtL5b//bEmkgNwA0C9m33m5Nnv1q
8ds2ZZ0tvwRos7YNdvxbPLt0X8eNDT+wNiJgOvAFm4PZInSPxyvQ/OO7IJDGDwr0mOcnTXApoII0
MVXoW+9uF99yMYd4AU+fVrmpkVr1iaQM1MxrgkD/loKzvUXeftNP9/mgSzuPwgvjd0iPZWAk1cGn
eJCUnXwJ1sCLZpT/GSNsbZjB6wq+v2E5GBZLhgNBdZAaxhf8VjfQT2IuZw0NEyZAdVjYdpXDvy2c
CuWDY0iRG9k/23SjGWm6Fdnvli6pITcwQ8u9M0yoCA+A8FwH+t3nHwXnhZ45ZvSiTUjkJzwN26jv
ju2Z7n9cHx0lNfJRmafQfAReZcFOTMgtkd6OJrkDS93AyWRQ0gWZVoCJDFIE9y2NTG/nMdbkmRtL
GpHG9bmgwMl2tHatUk0r1vr5qSVR8etqnC4EILJdrJyXaQEuCaf807KauF9uDX12bMao6aqe370U
hb0yNlt2xCLrJ8fwmTlukIvGiuducnx02+7ZWmvB7zhp0IJQ0iaWBGc+AvGIO9WeUtGDXfOQ0DAN
zR26xo1jshPBtohXCf7QeG3O43oMggcsqWI5hDiPr9UscEN0UqgkR7cHXin+125rLM3CYcj084vg
b6N2Xe2oCcJe2XUjRfFaTn0d1gxOY/KH6495PBoWhW35ETuSXteww0svR7IP7lXelQ7PSoZDd8F6
ausHzHKQDlDwx6FRafwscznpALzSZWWoQ/VHmN1PDsWQLOufiaCoThZcLViI5YnxYqWF2s0JMpTH
OquO7ls0t7VKj3qc++gdOrAeIlEKmST35e9/enqmL4s48Co1jMjt1ImZY8lLe6k/FXW7z3x8D4H4
HBqbdjXKZe4joNXH72jjkmQDC9hEUh+ezhPH+b5Ndkb08NxvCaYMTxpvXwbHiEakNlslJWXlCVqn
Fa+vWqXVEXMbMAxZbFe0ze40KqcpOfk8yKuikFt+4VWtyiGfB7hOkBsuXoKTCU7Y6B33VnHvigok
OoIyD2Ai0f35VPvhZUHlkijwc+MakwTqXN6mOHHopvVfkKpWKXSBx7gmXguBWPP3tJeMIsRwhfpo
U/2nwTuFJ389fFEKKDJdJBOpS+dW3TAqRwJLwM2QNA9IurfpSSPdLaXm7JSmVWypbosqhmPxQzQm
EFjZ0MF7820j4e1wH6zFOWAj803FsuaU13FUJcaW4LvoZG1qzCwzJ6qSaVlBaxUi7GTGqz03zS1z
gKfHEo0eIRQY1BmYta1ZWl8YzCe5MKiyJXymuH7Nr8eAL93tpcYqNChe0BHrqcnTF4hZ/i4C77XD
Ikc0xnE/WABRBKD0jKJ5A3tItmfVLpMzWNAbQETpt5zVLjc70WzSMUMyZuYriMgPsL0beH+X/oIg
g9x9W0lSniU/MiyLIzOpm33pWQ0ta+rOzD+ENhHDcJgNGjFpDoPk3Nzc0iV0z1b3wqWDimEMBmTL
SQ5DkqZjTe4HRNPSRookPG5yJo7kIY4W0F5b0Xfik5JxReOZDGneGYHcZa1tvinhz9vZt01tmZK0
e+dCAUIdRaZNhzZmUiqKVP7S/JccXpm9X7eRULm8wKeQfbDN/tS2JbEghCUiRTNGVUUAiWi446kx
FgbZewkS3h8J97ci+ifzsA4/hVjWPLKeJ9BWsiCqnuqCeqAcD/GUr0hQgW5z7tKaLfQgcnnzwSoo
tBzOjodUJN4AijAdedqAF+okG9O4ZWuvfRShEozByMPaRnzea6sC2eWtlohU42C/VJtYBVQoOQpK
ao/XxttZST8KK0a6ljHfDVqmDSYvgAEcqGwuo3ycyLqFgyHdtA2X+2q7PhxwBvajId9sBhddDdD/
vAY84sfFlmQ0ewlTEeGakCu3C6+TMVY6T6sWo2RF0tCph9qZaMEru3N0tKO8NZTj2rZz899eSd1c
0wFDlwgBXLmkq8jOxDyjNNw0JPvVyFGTR9afyMBYE3hCrqikaSAcWf82jBzWqvW8rxoz1N0f8P7v
if9Qq5OoHOqwP+MExu0xqlAGY5JZIpG3z6Wcjx/4i23RQXB9jXYp8Etm20kGKuk4Euhl/x0cSjNK
C5zXNQhHmx+5JNV1I7NuxniWJKszmVpQDplaz982vgDeSO8/UAFKe+tudXBQxwnqUEYQPbc5OoGc
EhksbkKukdjtiE/FkhIFFvyq2WpF83n2DX2/yALAHMqEuYn5Ym9wYD4Pf0gdkgBI/OQx9q0xq2gy
x6Rb3d/oIaaaWNkIbB6azGLE/UDEpTa8zBiKCZD01yywt47NmbdJa4Ik1e8W9nSPZgEN2Ln9rNdf
a/84PLRvmYMKW92leKXMITe6N2QmMvlp7AsioiQKA3cCqf7E6yj1y273EJlESBvgBGae3JmvNd0i
vtOugPV2HCLkTA4N/+WQ9vHo4/z48Vb0GFZP6WIwmLQco/aMJ/US3LOcOrpV8jKfxKGJBdxIC/Sz
6y+l56/kKzw6ymJqhppRMmzS7xvcfdwigsnYTnq/69ty0HHSQI+UCXAfcNObQ4CT7KpjbBWUXry5
zP/b281BZOpFI7pPCWH2kcb0C0L7Fo4PfY+AQkjhPtJm4+AejnrQaV2XT9pohWeH8PdlvEn413Vb
I+nJiOgCp2Xdr4HdTvmbzXEPdIKEJOBq70zerF54ZziuHe9A7jYWbTDqbIkoBw0u4rYq9bLwORQp
qg0j9tbEP7/nHpwb2Evza+luuDXoKR2pB2XgiVrLbbZ0O8imH/o8T9bg0V1XQtz7j57XC+zMSdZV
POO5S/MqSs6Iv9MQe9OJLt84PCcT/rS515vEAMcOpQm70u3wlnGP/MWITnSBi2+Vb0YMEOr57AZl
RPayabLqUuvd5pV21tT5djhGM2Sem6oNEAJg9ENRL4RGQ4bc8NxXKrXHYhi3q2GawZZbceiKhn1V
WNDvntFIQbJjUrn7KSoyuqJdrMKAm1l45uHhZQvjqL+4VQqoDQUYRbriFMY9p+KGlHMnBt/4+Nt8
LQooNW4ZSMejRNM3DUWwL7t0d9zuFCOfTRgqSECQghfooFo/AOGpgbXCFlaMrnzP4tuo2+WCE3Cb
cng3TjFHMuia/MJiUIlS4BK6kt29THkykYEQ1nZlOa44mQVzlm8JiFil8zXCxVCOiM/xmDcLFYlS
UbivNttq9IUXMY4fhpZmzVjaH79pkmqLyKVfj+KU0/DjykrgHiG3HN2egIcm4tbIp0tnKDGnyFBT
CU4EUw2OiddBtbFACejZ/dZQGoGhKUBVCKkdYj1w4XidzxQ6gbjZLsqAGwPl3NsRydu5xsZ/BbLP
5JHLI9EbpZGM8kgggpgAFN4fdaxi/5CoNPGlDs3doJcD+mNJGw3/jIGErGz4arxF735OHra/rp70
4ExaHerXYTXhVGv/DDBfzvacptIUq3vbxwIic5MXrUdVIPY2FkvgddPuNqUnnrdRhUvdiSWL+fv2
7TIDLLjVhp1QHMT6SIO0xlRl2g7ZAjJJw3tAESTvT/alEwxp/POCLkdos4EqMF56ENhW/gFvGuk8
SmPBqjQw7TbFU/Nty/zozQZNSn+VmL3KiWpTf9NnnI9CVGyZjRa17GY2fP2c2MehUBQqoAyQhwFN
VKeZzkw243nf4Bd1TlQC7EAzLLsLzDrf54fc2cwHYjOA/hwXd2ZORNOVu4WRt7ZA4QcZW+HdPwZP
4VWOUgEyDAShtuQrsiVFXYe2oikeCdesoY5Q+Vs+Nfw25RKUB9f+KqlemwHM1W4XlaMfKjEe9MIO
FovwqmAig0uwoumchgLmzipR6If0S2r4AQn5rUUrB7kMSBUNK5ViktaLsmRjueiIr4Mstf2hoRbR
juFOCxgn0zS99ABBLwpbhVslIp1/PdMVA14GJgGo3Okz+1T6pxHtnpIHAgdHzr+PLIMYRYQV25+h
2IrbP+8WvyJy900AKnrWGYjrOZdtSAF67VG8hMUL6WlHRWhD6ziUvzUQY4NhDHtQbu3oCh+xLR08
z0gXRdlVk9RDHx3zjwol0ebov/7zG7UG3sVAJGtqpQGAQfaHedT6cJvmIKvFNn9foFvvDMMK1eTf
+46qrPmhcsgqDkbBxsTSfZQdY3a3M4RuUXUVpzcloFl9Q9PsBu6asj9w41Pxcl+xqRnT4gHBoc/X
tyWfsC9aGTi7Uma48sq0T6FBDPpzCQSfpQh1PPaL29kO1JBPh7fBxRuXGu/uPfCZ3WGGeNeoibq0
AyGhdVfQobG79JPZWh2Ic/jJIjm11O3TpwuGHcZ0XaxkBPNHZB+rFW7+gljxk5jWbWTf0gj7d0gc
LWx6qmJt0SzfwxAz+BgNwWdC0B4IABS9w3nD5lEah3D+zPTlvGtbkx9hqzNi90UQghV0qnRp+3MV
XjFw6U5FPnPshuhn4hgJwNepJEhZN1i15gz7s+h1KbGNCENOo6+rKcbeEkNvuZMRh6dnaL4q8v0r
/bQygNU+zGjn0ZNx85QDa2c8FsTq4UOk8H3nt8FUd+o1/R5lsV/91GQBWCO8+MU3wrkbDj6QT7U6
3ADgvBis49EtUOK0cZQqqqMRSzCezk0fq7LN6fMIA5ByCrw1UU7Zv9IiQv/SvSotgA/wiT67Eruj
2vO6j3JeLABdM7KcQUm7gxGPl5PQVBDMXfXBuNjkZSNcXcXgT6lT8ib+Ceuc7qzNfWditunsGtb4
+goSx9n4hw6nbD8npLgolcaqwopp0Y4r6Vy/PTedhiFgv5izIca2qnBEeoIeXhVqyhNl+dvTwwcX
hql2v3hVPyFnl7eP/rY0qzTzPaveD9yFNH2sgSK6v3K3qJ7JD2A1GwFoev1HQQndCWP+7G3QslBF
OJWwteO/qg7uCWmek9CnxLtGmfogle1mAQsIjDSrkao6ssIvtsLkXhV+8RMyEHaZe55yWx0TiXg3
9NEUF4I8B51NPii+lOQPQytvYYTSVisLbqxCcO+OBbYuTGtyJIhMaSSSHL8Q2mbSfdenJ5n9HZAb
WnnILjxKW9BZaf71qz02STbz+CykILKAGPvh9p32PR2bM5SxXt8WnWPo//3njwkwx5ib1kJEXP7X
vik1VlGsSy71wiIIMopD+y3JIJEYDnczDrDJJM5BYBlESnqGteApVRqh8jZz2tuoZwdLKDZs7uZt
To0YsqLyBTALVJJM+okrqrntWItTORtvpVLpOFnwPeRk66ddSWOzLgXC0B50FBTm6xmla4lkZISU
7tu+9JF4EaLmDSw/IDBM7adKJn4aDS9JwrC9ypnei2RmxVTPw0cM0g2rU13zpXul4e4BQNcQfON1
jOfgdotL00gMh0DJPcDoAcsAKEdLpTr6QUbL357dr43BZbs7slEGK6Ke0jkqsB7PRKyrJwnYXBja
4MbUcSyzkr+sQLaec1oCtV8efNIZHF5k4BPd6xbhjiGiS4hnfbNXskMrxV6R5N5sImF518BB0NQC
WADRO96lihl6LvNU/wOHxoc3jNwAcU4mxJ9SuyuabKpRZJEDTLJw06+5INTdwksAtccFNWJdqnCj
oPzmTBdhPmFBKauVe+vWPF4fVHhwH8LKS/Y4BawQjen/VKuH9jfVHCNsMlprrYPHp5Ng/wKLB0c2
CCUfjJy8N23eithAmpPMQjbFDNgsiMP8gtreFOb34OpjQmNASOTcc1MscU53g9n4iS76+FyRF6iT
ttQF5t4SsiyqP08jAsinIdreO2mvT07sz1JG10QXIk0jW/oCZvSz314worB1+XtwPleYD7aGHl/X
14l/lJuQh4EfKNd5q+U0HB+WN5cRJa2cy1GiBLy6doybQtzh7DZPfcIq6+Dfw0vCrACR9cU29qYB
6L0/lDtZiE7ntML5rQiFdogi9EsvdYDWPfzSxgzOjJgEXjIzUewNsZwY0BzMF8Rc9lGYhYY+WO2l
ouJcuKcFgsh148lpgmBYrdb9M8PsDZUbdqpOMWS3RXU4RtF0KWKUFmW1QK7n6KXPAa+3aXbzBqCW
/1CtQ9aHUkO/Hixo2CUxq7D8Scki22M+Fd3fapof2F3CTauBggr2QWUAbShR1GfGtgDP5x2m7Eoz
Gk+9psL8FnOm6EttcnOi2YScW0BiV7vEef+W/NjCQ8WADHXhkug/tISVldVth5QwJtsUb568bqd+
Fgh5+HtXEEDMfibMG7lmfZAF213N8usRMQGEfoW/mS8pL1u8O7hmK0Jb4t+9bj7D/RH0td24Aqeh
MSfdVMG+94H0cK6Ibm4CTcVV/5QSPtCBBU+Ogdk9buiuda3j6k8eCudH7LW54Fxi2BO1R1bHwK9G
q0+yNi2BKRN760ItzFjBV6N9YfKC1nwjvAERdBxvgQWnkmswXC4So4FjwqNVIgUQzHXrbkT8xRjP
1HSdWBek0wK7Dk6CRd0HEKNS59Qcp7CzjThB402eR4MYfGteGjW6lkSddCcJbImgkNDL8RFLOSqq
ZU6a3xyUNtffyRjJ3FXcUwt6Opu+hYrzH3KIP2vR0ZyXkIAuAv8/HmxF9LU6/h6PMGAwU3dap1wl
fvyqa15pbL0l+0XGqyS4MQrlnUCsl1JscoTHIwGba3LCI7VkY60mh/k5hg1NjXGCs3XoSXJji/IY
tPp1qAlyqz4RYlm2/g/HpN4Y9KONn2LTV4OmhAaI2HWEDJTrHJy1zMvARvasoKOVlb4/uWu1ptiY
6jpOCLuqK67v+rQep4QZS6U4VCsg+TXFRqdJVrQHle3QYq6ZDyVQMq8FUJnLxmkKdWd/geZwhu2q
wrhKDsQSAgsVDN2kiPqlnqdQU9gPpo90D7nAgckBnDjfrjn/YKzCKH7AGhS6w+KQrpaL5DmjaDff
tSbi2OdCxV9GI6JZN0Xgx6brPCpKzRcvFgfHErm433jcwLMMYtoE3C05M55jT8/Uf209gCOmuSDH
e1f2qVB8XtJxYwQlX9OyWzCjCfd1et7rUwDZbU1lwasNpx8GJT82OlleKlyJv+5Do49seku3SbvZ
Qdpo73gIw9o3aangWkcgXvFZ/CvFIgyF/YwkgBjbAtBU3OfQ9a5pTvPNP5WEcmNlwLHf0RB+7Uf5
85aueh647+Ybv6NsBfUea4yu97xhTlV75EwaJwM4Coex2KFF6AeqN9MPEwGj/W8cGUsL5Mfhx3YV
5S1JC6PPDe+B8a466K/6avVuqRxkVTb2KB2UUpVT5yHSptZBBM78qcRzHyeiXcb3z9welYduv+3m
p8YdBGRAcZK3miTJFYUg7cDdfI4QJPuuhZqGDGYwaQLV9Sh5s9jej+NI8g13x8piS8MSlsansgBH
3s9CxCp7lAD0WcOVSse/cjWjFz0pq72/Ooh0e6SJ+zsKw1+aHn4+l4lpTOu1ch156ZfoUY8npwCg
kQ9rcPi7vXkArZHneJ3zm7s+/dZPlkNc4hSFtnWTHgPt+/pNIAkGUDuH5cq9wo7/nsdX2EPUNJJz
P0Zlf+qvOIj+A3wZKc0ph3PwtbXxOKQBn+iUpGaoiZAhnnT4I3CzYmwl2Ii8D96K2OOnLruXxB/5
DoEbNBGox3sNtV1HRh8mty8kONPimfywukxUGcdKvKtMcgM3z6vwhpLevTUcImlTH2DjGT38l+jn
OdQBBe+bNAKELp3gFJMfkTrRy0wNqoJF0vsncgWJjuI/T1/F4g8sOCdIE4Sj1dj9g4SipaDZ2di6
WHA+SKheo/QczGyot1Qu1DexM7zrBRyIodCn10aByJPbw65p/FtAyMU7re8lyfuPONO5Vo9LQpZ2
UTloZVVfW3O0ndjEGtvH3x25krVPyr7Mc5dHG5gjtl0smdqUe8nndVCnpX85niHJCAoRm869wi+G
FpcaQHKie0B0yzMNZvw2mAARPWa9tTvNG14jBbjFZbtVfg6Ek2r6rLN7fP2EE/DzCYz5OHpAUxCY
SUQs1kJcA6GEZYoYrY2Otrm2SYOjqmUSOSr5RmqRZIuI0al8DkP/VAMX48+qKtfhJ+mQNqovk6gD
CfwSy2e81DoDZwKSX7003rHHyBXZADb/4tMpjTyNRUU/HkHqly6l1xCfROhACrJ4pm/P1/KU/NzN
s4If5VrqgBSzZTF7pX4e0Xlnfa4IzRpJBQG4NrH/y1avZIhG9q4PidbWTPPhIPS0rUdJM7ZB/VDv
SoUu0qfishP41rdCpkvDFRYkbCml7ws1Ai4hKhAQxvGwXDNbaF+bgc6+xEr8HQJuZBxHBMkG3ITz
kunI3XJT2EF5jagO4J8VMFoC7h2WY2m87Vgou4De3BhaExnLz5Mp+Ito1t5zTF+pp2ug1onjPisJ
f88Ff0Ex/X7StxUPs+JLPkcNdUBspyHx0XE/W2ql3KYov2b0hIpKab+7aHTjZ2aN6jSnM56Te7W3
a6X8gKo+MvaPnvyuatsUdZ17x0c9GSTqUAtkQxHbo/DF0NOI5F79mwogiYpPawwBQbm0I+fPvsQm
bpcpZdO0vRkAkdzO/Q+5QJO4fSpiiUug918CFFg32Oy6mBXz1Q+Pw8MJkridbvBuagbV4i5cXHHJ
VRGGUxSg+yrloOWvPvwkt/lrdYtyi/LJSV/SEtG/iIGp3/sEaA28ENqe8F/zP2ciEc0FEdtta1Nw
HGBx+k/mteau/sDoHL+tUnZKnY3v5fKkKFpXXfdftAld5lbINcSsUZwQM2n13EKbsFClrevs8HuC
sH4xv0WqhehuvcTjAYfYj3J/EjBnPqaSX5BedndKVh9ruNzMASJfn4/CbNBxp18gNDLRgcAz2Cqx
hHdle7qx4vTRoMo7Lta16+wodpY7lOVc8C/GOcFWQ38BEt9xidK48866kEtvxQ/Y3VS4quQuZByz
4HM+trWbVVjMc0W/wv1R53iWqyqCZx+2TiILGoNQDy//U8zu8feZBd3A1j4ickVQTwgRsc4BAN7e
C8wjVSbgPtdp2LJYIXZh+OBwHQNeLcaUuhAqQYggqcsR8NgpHw+IlvVb6dOpHljRe2jETEMacHHY
EhavzUEUTt8BMyLc/OjMMp/53AkIZOyJx9GVsU7JJhTAT792coqCfpW8N88nNwdhtcHcac7loMS2
RBX8FZR3BrvWrDo4EM8GjrnfDrputCqGZNd5QUCxiyt4bMRWbjQBWSs8ASZQbjhAhtWXxc3Ds9+N
lpW9mKwxd0qfam3LlZrzEsB61OOcJ2LUqZ6n8sot2mAkuHAFtzd82EmOx4mSlrj7mVH2Sm5Mr377
wSZK41dYtaUVmdKbheb8hztUV2IXJiEcj4FIJGaAGKcKKDeJ7+r6A122yiLv3cV0PH1ZsT9WIdQD
uJqWpFAtYayZmRw5ErEenb2BVlR21C87TR+/V25ufCsmveUr3KZc3EtpwXYdu/5saZu31d/MiCWL
evUEcIU6EszW5H1y68TGY3DdYK3qcYlBUeHZ6Lk7QTNVntCDQohMxku2sVpenMrMmuLo8T6K4UAx
r3rF118xBC8OIRNXKJnN/VwERqv0d9ALi0aV5VbEFZnNg3YkWWM8MW9/qUFLNp+69SXqoO/Xl3AK
Bdj62UGuCN2xz229i0aD3LcWQaKi3M5ybu1t5ipeVZdE2nL3Ok1t/+JmWHleVYQoRVLHYe/8zV6Z
FMtvAbvI6CXW6GNDRirkqPpXnKh5HfIFecd4bRex6rGNl30fc1xtl3/CIS0qf3bLVZ5lqthjmQza
lnxd5bHATi63ZAuKqOTF+YNfydOrQdo/eXdmegemaCRNImGHe91ic2baG7jZjjyjA20xLKr9Q6hE
oRYUEzmsI5zTRa/ZYh2Uy8hJfb7Asr6m5ZF/WKy/I0fLsdsShWPuU00LXpEZCefmhRcIRaYGk9Ig
iMx0LR1eqcfin2X4t4troKkMhQlQ73/pPCgOMhdClNGKnftADtFkini+1iOco+Y6f6mUeyBLt33Q
DVVP13EWMT9NXFC4cwrFIiu2mORYmxIBiCtzNgCpV6mjefT+1HpuAEDqgvCjY3pOJKpPbN86eQdh
Rn2mB438paxwYrBmhTcAkT71xP7ZUsoIKq1yAQ+yJ/IN3TrvKbAe2/tBAs1tg7vwgfuCdZInVtMv
qwb8+DNI0gOErf12GFjW+xH1uTNfE+72QrxFu6CkLVGwn0Mnmp7UM4gRRN/HWprYpdM/jQt3xQK1
F5wZBF4y+ZG7lE06oFfk6Hw/ImKtFeN6KotZFoHltBmCweMpbjE6m73DwFNHCqDTus9fqtrYgPCV
FA2rhsjy0bDVqVviaxqOtcIuFlBOR8vMoARwJuEXMiXvb9+ESrPLn9TS3EhVYTH8o6HdaP42eaTh
FvKHwv5ciZkiDDFlFTx3ctmk2uij9TOwvx90Lv+NPMDuKHvijH8qnuaK7+m83SvucU0ejY72unsj
jxOR05iY5bZxWvQXbvdTJjcZa5Nkrs7sITyJusdmIGsUcIjF2h+5Ysnnydv5SjUdyKg9xKu8tR18
t6zQ7XGY/k3dJuAFWj4/5yKExLm8P/+hJSIAoZ7RGmrMXnZ3QBomDnfDa6vzddi7KNehMVZ/k37E
ry1OHc7X9GsD5qZTgMDYtclRC4e89zj/tnVXp0ur8iqR+TkyMNiNYhWm9MEZ+1DHz2L0anzXM/V0
zSmsXKh2oSnUY8mOOTyJsvNFT+K4Cmjp6ndm6bWgbFBmAjzOfEpq6momimR2M1lRGap3TtrGgRfw
XrufpMj0jcUx6jgeEbLlfk2fj2GHzJCji3LyQYatweNRLHP47YaZ7MP7080XFVLYlzN/4XdQjJof
xbKkOtgW+0I2qLhuTESAoGXTFE3zuVPb72pwtNx6d1oqAJYn3527KjbjIbyDKO5aLBlqEqI7L/na
0OaFWu/vojAYpA088NLQv3n2oXky6CsgOkxTth13jll3kEM0HV0N50fABKgcshbB4gOH6AnVxT0L
+VtHDDozBniC4NXaV2HzLiHYS+OhA1H/uF5bdh6ibYKL2GO5TnBPJovB8bSf5cr/Ka18UWqwokse
HDszr+BHyJ/ZVmiNJTHGcW3jbqujBdjbKsuqvWzFX0fUsubBcoz8BggBlQ25xMNdS8wo+o0BkbG3
NiPkddITx8UKYijRw76DA78b4d0sdq1LK1DYNlbZ39OhlITmqmefvcrw7fAtnnCYVeuFAv0iqPRe
aiHfK/kUBWmgmg5xMJ0MVJlEDeXnYOEQ04dh3e2Yp8YXMZtsNREL3lcuHhSu52+MonJSanfBnYJV
rXVY376NTtAb7l2RzDE+rjd8UqVdLYarcYB7cRCf3V9Vr2UzEGKpiRj1lZFazN9rYV/Opeg1AmOb
bV0D2MmG2JGIzjGVLDo9yr69MdZvqYMXK5DviUxV2j5F3zTS9vDUJrtwHuGdRJbfisd36z0FWE4d
+ZXoRfT0xMuzyDvdbaWOe2D3BkVgMJd97tF8lQHKaswjF5ssn436dprAIgh8q5OLToMO2gEcM0jP
5VQAxngvg35d1zX/shE1v8zIRI/WkrYGDVX70XOJFgpM8Z6oopTl6qcW3/jA8du4W1112+EsHIKi
6x1g6xmO3xFN2OKymAggdowtURcwYxqdxjEeu6/I1XFgVJg+KT99uyc8oRiRuhrVE+nL48hFqIiu
xoBFU721Wzc3rTEJj0jdMd/LHUm/t51nK373aHpwVZkpF7FZPkrTAIsektzZpLDJlsguSEMVvzXi
OAUUKm96Lu46B+gqkEoxliIAdnfHrqY9HSz4k4hNLWvHy53+ZrXryDBHAL32IbSaGTqOVSNQ/t1X
qEeOEC3+c6CARFOUlY+eIdeQBRRsrm2bRYhVNqBVGS4yT/7NudviVjxi4L+bI8nCDPB78XcvbINp
LVcP8bN33pb/E7EBJ9OOu3hoviNYA5oOf7RmYTrUsaPQvHc72vOzP+IpVkAFEfMIuVSgkA0QBuKd
/Bp4xi4yfcRnCut887TjWEFhtT6dKbbzs3Nq6tQjQ+zeJrKFg3XSNc1kheiTgw0j/N60R62yIUsI
n3pT6Q98qOw4LMXcA5GkeqNVqWO/7/9LwlpjVGH9M62XL3DnnZlTEXNEeNqpYQV5egGhZY8z1b7h
pG+OzlSGrbC5MY9HmBfYyGTOeoYvPAHfayPAtUKKIuGQthsZ3dgw/SEk0WTzLuMWTRWyQGmCxfOn
zFKrFz5Bd6Wx0D6J1ZW4kirx5AXRD4r65LWs8YH8gGCEql7V5uHxOl4iEzK02OFyTHjgZjfw16FL
ZCzGBznr/ohAAbJK/wbz49B88ybEzll0DM6Ij9RKXCQjDHi8+mw79zWWHx+5uHnUGW4HFtiDtfM2
/KIJvzATjLlceDrey2C6N4LY/Yp4Nt1kWgXBw6Hl43tmXZkVAdkFLWNC4TWBkUTozTchLuo2Wx34
BCRNn+ozqBIy+F9waGQ7Vk1xB0RxrrAskOQLCoKYcFloyYk6pVOUvSuiAXNPi/9fOc9Bfcgf1YcF
UPvBsdUwWjWHaQjClEtgZDFJuVtTcQAz7z7SjkJT8QGGKMTe+Q1qtilJ445YgIa3uBgOKI0dwrz8
QZ0yKwJifm15s9fl2zw1z2c10JKRk6DBh2XorfeszpuMUDuuCrOs7iizbAaAyXzEXj8El4E/t+IE
GCpbr4JSIi5OU/cmYczoZGSdT8vlt4q+xX0je8BcNI4rv2H8ThNwG3h3wpatFJog6AOyiM9G5TeI
/OSPCmWcn289gw7btwN3vPK5XPqAMm1KYBjCDRXsFFAGDEVCsLIOxYQxL6I3fOWgjaTKgw9bVunq
OxUtfZCcVON/GNk2heqppZfrekjJJ9M/5YL+Gjqol0Gb7nCNhzZa81B604OeRrTAmqPkt8fn4nZD
QLw3NQC5UxMaMKk8wYi3Zju3yNz83xYQ182cidv5U1byWn7jIFcVG8CSYdaE5RLhr61GpUKVzIlm
Te6G/6ZONGepIfrRjCPJlVqNIwK93+KGQhrUNyzo7kC0ZyVK8flhNKLOlTw8Shx451S0J4z3F+qj
eSNFFvLe2FSqsQnCkz9RgzBlbhlPFatucOJD9bdW4p75zU2+1SoopOMpfIOufTkUUaLlan6nIfkN
tEmx6B51k0deBOE5IDagKYNm4IBQqVo4PQWOiUzno3vFaEOskCcJP+vsiSScbKO+G59b3wurfcZR
7vZAvCHZSNCQng+9Qu/30XFaxkoMJY774pVZ3rAUO5ZWId6d/y/OqwibMgKtppXRPt3JEpIw8VgK
+mtpjqpCjgYEbVH2QfbuZ+bIdzZPPyVq8uTMEXGDt+wIpPSQgHsnq2NozqpsSCcW+MO+YBISjJnp
rtjTL+3SSXsQHSQcqr3s4wSMBxomZlnArSOW9Q36WxX4gYA6MVdGEnWQYyUOVGXeszMGc0Q2hY1J
hpWFM3Y0091G7NKehVKk1tzYUogGUruSxjWBU7/Ge5b+5Lktiyhp1WY4kDL05oC1itotLWmo+KeL
XWTDEgHQ9TJStwEgBaPuJjtMp2fe3X3f4LoAuyMwItBUzVUFuiQ57Aw/2Yz22ZbZhXwAcefSDj0t
rQmDgbVAkiuIYiTb/80v3tjBbvXyZmQrd8vPPApsZ+4bz3yk0yRqXjiu4K0nIPZlG1JDq1QabXS9
NdjROuAbh+UnYQgZTGolqEM+uBBO4sHS+A0tzr5zst1Qyrn/4K6YSWKdp9A1AtyJjWoA3k92fEmi
vQDgBp6cioRqbdt1yslcxqx3NSKwDS+1iJxgBHyy2AgsIe+DswMMGIy5aTMntnGnzReSlpJOYeo0
1FMt8YDGuZ06WVNsAenNfH7lNze99mOWFCAnEykMnYvYO5pYyw3uurJnDmgSMlcXYQ/pMsMqfSWp
NCSYzXHNhwkswSeUSMQKZQYpcVAmM9riLDzAf5TXVSywdkht/Tq/coJ61ze/5GVipBdx8/vBOXIZ
LuKp2KmF/eysI1M277rqcPlaGdU7gzuWd/bvbRLXdcvV9VLx+rb9qLpPVdqbWY5Ac6FDtmomoBV0
XruXBltbycN4VQ9MhQ21rT2U+7TL8EEiAe5QJJ8GSJ30B66sB+GmNb45sbUNfFIp8mxLOeaetQfh
OPgbDPseClOmvuSfjER3EmtwV4Rc10sQ1VH38o4eLnHWWbLrtRg1UTWj7wtXy3qrKjbUNAl9Es5L
XKkLV5Fnfc1vzl0K7M1lQwyjiDZDy0bjvAkt0D/r9hPWCVFc6j0DdmvVJTMmdh0T80UGJZ19uDvQ
LyTyXTNggOMrP3tice2kjPFAahD8SKNr5iMiglr4Tf91dzssBIMosmXKQkzhsBJ2/1kYX9hyPGt0
OZA+Sicc8X0RTGvFQ4UPC2kOEqUqSnPaZ5Sx+3/3ECAekQ4OK8gaO5FQI5KjP3fS1UQYFDkJ2Y2s
V9g1ZKyN0/dH0x3NfNat01R44zjTebrnuiBNhA9slMuCmOXPKu2k75tnJvwRGA7GIf6iUI/wl+VX
VH0izJB8+dVilHLBQRtISFIe1w7wkB15toHxHUrEk5YQZc+0ihe/vcwp8FIgU5D4sdNMdZrulPAl
VRgGuBOOQhrOtwapd1qLwwrcGM1OLj0ntM2OeCdLWUdVxJGIqyGoC9CDwsv+FcLVYJ4F70tpJro/
4gp5/fudIZB8y4fMMw8Y5sq3spmXe0gK0YsSirRCxIAI3DOXEeP2DTIk546lnhsrijg/HaCZOY6j
dbmp5sO0jV7KAo3T/AcNf+LMP/0E8uowHZzLG6FOpRgvdafXx+4h9eQ34Dh39q9ELbPyOKRyCK2u
MgTvHH6Wa0pfdl8Vg8R6mYVo012zIR68Jg9mI3ZlFi0WLjNX1ZdfJID/V8jXFdSFgMRdaejEspqx
phMItA6Ej++gjjSnyMMPAh7FknREq9hN0wkbZI0EDNuTGiXME8wjZpcLX/ofqNz+cNXAZBa0yMRJ
LnrJjLXhAFZ9zOiU/2RXxIjU7KgWd298KTTJCjShTqFGJTu3aoKLgMZ3Lxq4I/c0cx+Fw64dckjC
ld+TWh4C3AR3PFnOD3rcIo/CbCHpEIsgd8uF+RwN0ojN5nwdkGRV7joNpqVCVWYVhtcSusXbgspx
9b6zvHt3k2vIimLVoaIhRw+P4vHVHg0RRxM1SlJRx5J1hrVrBdZq48+TEauaSY8YlRtfRpQupEvh
G+VdNlFhemitBaGN0q3Ld4mXI/RR8UMWmwTOevlJJ5Q8xlguSOOxkNdK+WSdZvx7aZqdc59QI0DX
IgdYdZRTtFCFkNXrV/yAgih0ZMll3wso+kpCX99slBrEaC0w5Jq6Mu+UW6MnVLdP7eL3gQEyCNHU
8HS8YHkkhaBtaXKN+e+JrBUCengszjD6pgXboRkiaT1EheMs6bCZGVXgFvpNNm8qpi13hyi+xWbG
kcCpIUW47KB/P0hDDjM5OU8zSD31qZy7X2BPQklm129S5m3bFmPNm3ncdF9gZ+spVxh9XcItT+Wo
pZgzhGpmjN/+jqUhiQnRuzXFXw4ESeYdXyfC8Gz/KTtgJAoZsr89YYJRTp+eF7b9yRE7r1H+NU1B
W55knygOLx14SSNrWAPXOrzpWJlRgJeAU0rhN2OYV/6Km6BTmk+GyUDlAPBQhbI618nktulC2aLt
qXh0wkieeDg3HP2OOfwUF4iqd4PCFW0SWcTO1zeYB8xe62L44RtkaAwEvBPRLy167htoe3mDWIth
cECt51Tj2yHH4CaRFD2W1NY4P1kBiy2jSE0WZrW27Op3hOlELXVbSQQE7C9rVUUi3dEDfulNn1FO
FCB1fEaRjA3h6JFeOCxRIQen+y8gMDVrbK9ixPy6fSxGLo9o7JDfAUsgV75iSAvPIV2L0MVd45AZ
MFrU1c9LHZbj0BlcU/JzET1BEspR5R7PR6TdT7oKSehF+Fln0kd8cn+PD9AYJSCjJ7ByFU1Qfkmi
Xd/LHpyPxS/GiiFioowkksy9b4krxJtVf2N6GsTf7INh/YRf3SV7Ulr4f5DqqSqh6GQy2JsbmQcH
izQTeHrp+ncnVJ6ecmBbcdj6/7yu6hL/ypx+VDbq328Jwk2Bp+h0HhZTewPkspHnXRfWz+joYkpc
wnp3CGbCk4e1WtsA8BiabtQTj/Rh7XmRM8YAmFXxf2RonuEzLt+hKt9XRmhscRPl1csRwEejsE4l
D/lAGCUcbiWFmSXuDUhws49Mk2CRQd1JsLZYNR1wvhRgEAfNMu2X6r6zezqaYcgTJZyYHhoS2b/I
FFdOQPcGaDUtdMqSLowMI/l8mh8+uDVYmEmyQREf3ZPxstODVq0nHYj/8oJUS9SNMCrGPNer2jxU
LHrWLTE6Udbb7kKMYlKyhizi63QM46MDHGYziRoz/nBQsiwKvzEle8FhP7exfWtpIAKgwBRnF2I0
WW59Jy+SQC5s9X4FB+kQA2fZM0EjHvVFCz+b/Jb4M80lcE9XO4q+aP/yjClAkzhlGCXwnPus1Y/D
mLZx2kbOnwewljmKTeUifmM6E2N6i/t7O+S/xAx4is5PbW4wOKAxGf2hieYIS+paztbOT2r270/z
Q1CD/irfkZb5jGkPMfG0Yy7Cxk/+N70AuSJ+c28jwlaBciw7LHHE78CHU8FNa4BygkIxCYMv8h62
E6r0dCMObNpzrte8w3w5IwWhFaGsk1C1hxWMlWQGQBPpmCUAuFCN2KEMJ1ElhbAnj668zSTIO+F7
qZMKfPaZpG9G8csRcpVGeCEbKzUz1gxpPPAO6BjnAeoznn6t6yHK0yxgTXS1DgMqL8Uo87pFav6i
X4g07g6Ilnj/JbnEjkn7Qs+1o0mLtYd0lw==
`protect end_protected
