`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QOjT/s4LGWTUmMFXwsJA2pMMxPr2D4/XXdjhv0LJP+skeP5lQH2lvU2aSpwKAJ8jhlp8MCDexr+e
UkiA2h07rg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XyX8/Ug5+Nl1VZuVZGqlYaBHBNUWmyO7QqBJnYAk0w7RomiX2+2FW9qf9sWFPV9rwtLYYU+It8O8
AsRjPz05XlZRIPlMtJ1ydUaSTXT8QQA+ZBE9SeCFMvcoFW0nHy2HmdaNXSEO2HBiplECZakfQ6aG
f/UC4u9BN1eVLbsiT8A=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
0AI57RnIf6/3DMSlMdq3dnyBcxkFKKPa1zJ501sWolVLvtH9XIL2dWWv5vm35gSVmL3vvxqZ1XRD
v150YgzEog1U9tHlJ2uKUbZI7uwx8jNpqJ7/cVttaIXuyH3dlyzIVOL0NTyMSRktgBTmba8VEwPm
acDcnAQd/DwBq16aDAg=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fRPh6hfnFJWoRbVSl8vPcQ4w8/+DxrnJMuR7QfpyusVtyK/p+JMMfYcA3lLg5DidTbJSY/UiuTj5
S3QlQUh3Th2OkmPoSCgVVZHNDll+QOMMpiv/3rIYKz7Vgl94/4ZNWH2iDZ6bJzIdPjcVoFJJ7nLl
W9BASh92MPxNG9IuRj3+zuzcYCqqbcE0lyoA4DWa+JZ8gYdiR+2Rb1brXEZCFr77GJ0XNlAOdngY
AA+dFy+TgkSw4hmuNXIw/KVvArVUQGPtvSSehnP7klnzDlsmvXxxHjN+EsEDe1Z1jqeY3fgkfZyY
1zcSuV52N32GJJK89/KsM/cIEW2t7+V3qR63+w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fmmki/A5lXpj56EAhjsdewolmWataCdDTkjztl3WzSxca5ucstuLUi93/7uukRmK+uRKQsECuo8e
ZnvMS+Oj+TsWScy+otx0IqEd3rxC2Q1YxXZP9RgMBWP2ILiBy2QpDQXWkJgc8P5Em9vC9rVOXvgP
F00dhZambETaYt3rf2MimyQqnfXHpaTcvXW3G+4UkzRgKfL9PVXxR0mTLm7Xn2jUda6r+wl+JRFU
epuhe5j+0e4ut09tZ57Sb6Ch6+5NxRfERWsiYPE+5KpCw4mXUFmoAVCnJd/BSyOsZWzFT/Rkyxcj
TFFaVcbWBpkAv/Q2iY4VYx4Av8PxH2GI1Oxbtg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sJ2EQuV3SJhywYiUGcaWCQBbFz4uh3NfFL9k6EmpvrneHMa/zg5d7zXzjhu2grzJrj7uPvqMFR9k
bujYt7RVRWFKQKuvmarWY7No7DKdZwKZLpMKW3N8cMFHNeIzfC7HlpUf05anS2i1vdoS7ToBD79b
HaTM9gLOC32Sca9Bf4wtF47/6NN2Gp3B8ruJSYodCtFrPPrK5x07V3fZfypWzMf/xoH73d7YX8hj
nEzw4+YaTYMdW1qdNTsu39200YQ9kq95GOR7g8dt70zE1JcrLcJoQ6LwaG4DYh5u8BrQFHZYjvUb
VwcIaCu8zw/zma4QIsVMwDl82hSh6EYahRR+OA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 175296)
`protect data_block
5EQjjrw+vidbEvJYB69q+QEv8BTTd1aHpnC5eBHc/1zOWFwFOHfiLDb9mEYwcURqEdGXh3oRNjH+
iYtAmdqMdU1l2zmO5JD/T4nPOSFghP8uHNibbmUDqrVeRJbMU0TKmQPE7AlVC/MLUKOMYkI3rrSd
93qN1WWwmEHxmhfRT2iL3yWVJrAd8rweT0ac2kVc8xgt4heLVH0tj8k1mvUvwv4IdoCxhhaGKNFY
Y0TtVVDyKSN+gRAMPa0+0w44Lr4tp7GLsxTmKIE2rPhaa84h7pf+mEOpzmnhFs0PZTajI336CduJ
s28tBtmCjIMH+VdYJBPrq77Ml21K5GynwtsXBA7cSnLmOKHZ0cb2lLak0Exym+d+VG/BjejHJI7c
2m4i9F0w8ijzQG8AlUiLSzgxMpNiZpirR37znhMvNjNTeQwO7vEQdnd6lv65pGEAKgJtpgzYVddP
XK8r5N0tx67iJsafByS3aC2wAAlNbfn5htrmjLuVlHOmEMsmaLH0DkZPTj+QgQ2fVlhGpEsdAapw
j+6tF1eo9MLUIOorGqoONG0FduzOfq2j3AWKM+UTujXLQtpt+RYMQ0Mhj8MgJW13GY1H1zMCyU3w
I+rZ/TQ8PJoqSds/3ar3oz7mwZxIeAvAhfkIWTW9IKHcnA/DgsDu0kBvvLzaDSCfi1TzdLkEyPPE
Xg96CY+HLCjLbmHrKf7jZ15YxeG3I7FlbskKYwq8Gy6CNcDh6PmOil1BD5W4o/Y/A7o3dEqXnla2
cS5HYIj6bLvrqydo7osjoeoKj6plXbeKv5xjua83cKueeV77giBi/vyXZKS+fh3HhkDeFiDfd1o6
ugn/lzwm25/xqn+TtncwGgrRs6aD0GEWK1u4W5HCpTfXZ4R1OPvklozdBr49KElKMnLyUDv6WCIF
6YYmPcbcEBjskdEoqQqUCupKVayZjLHEtV0OGgER9MeFGAZi21adSOzfNnFSumDXflFH/IwbctW1
mOYczTX8ngXbQIprEVb36jxSheOFutsO2jo5+VKDURmbBaMBGlBkmRYxKg8Bx/oFsRyXrARV/MfO
dMjWNDW/HDhgLLV8YMcVPqZU0QhGOiIJR59XX4Y1BORp/3F5PNxjNIe/pKoqjNfeWAqnfgk81Jhe
27gjbeez52dQIBHixNji6bGD9aJv44x2vrBT+W1kCir8VM5PKHZBsqT+7CXW1TvbEnaQ3+hAf9Tz
azcZhBLAEvR1KYZTYam6tGQpxAENLOWlQUJl9B1DxgE/KGuEm5Z8n2N8vK7rx5rqWknGxjfKRrvp
fLZ9roOAkkhuirkCPzLDL+Le/8Xlsn/pcqsU6gNTgrdQEOLIDs/c/E1msUT4vqcCPc1sfCYXv1zi
TB+zDjdost4zTf8/XGvC6Ijkx2BP7XBca2LjXpK94ScbEQYOG8hFqi8RWLCgm/V8VigZwDX+jvNf
1pPI4BVhEvzxjRQcNvDCSyyQqbRJAmUzAZIONqOhhYOhSWLuZM3iEaYHIafEb2amqjRJ/YPHktzf
1DSbURc0FcMQqu98SfDYCcOiCFrAY/wb2SR9Cd6CuQylkawzA2aDJTABXGAEv3j+UrcGWqHvFFq0
8LnSECQfAMYidNGiFArG7Ye1CMs835taQQw2pBa1UeeWR/E3O89MLV9phLk2B2mlPPp6GEZ8fm8B
YmTKf6FCKHxssRqJV2DPhzuKJVdL3Y2h4nUdHIqSB4Rx1XaR7+KFHEwepd7I/9mmiTnyvqd2ofkV
Ic9t60xr+LYXvCdjWpTx+Nqx4pXb79Fg9auIKxM+YVuU0acwAEGDWkjpirVZfdNAjNyfbR9mdcMH
8hcle3j9xw3RVaB4TnMQpcN2QC8whi8GvZ1pKJgXMZ9PlLOL8PENBysfxcGZfhTjcSjPj/qspVuP
I9AnEQNozKyK64yuqNwteD4c2Y7tiOnuaBDBSGD7TJSFyfvUzRPxqo54xgY6CTukoLVHTfO88FFu
xi3uNHSkxXx76LsAag2W29Rmr0BCwpbGbbWHqwlgyvbzSCELgQOm6a9U8C2yK//CuuLEgu0JKzwc
0344YIbe/CAxyHvWq4bqNFF5ccwpxfBNJzTNWB8kojS55A+NbcSCCcuiFXngGEGzgrPsBD+GX9mD
K7IAWkLI4u0U6D/MMxWvasEgpzhB0uZcN10DBxYrjsLsbN3yyxfIlZF7e1dwDBPE6Y6DvQYZv90a
haetT8XTHqxWPZCJmtVxJWbdrCG/tpyB19AlaebmMGxyEqQQsZW+d6uEqOAbacNdUOOyWp2jVOdi
6oHv55QS7SZ4/mY18UCh+3BQCRVOHlCD76glr04lVGFFYyUPF98fIqZ/eobR5kKdWXgNo4+YC/JW
JdAKBNSEqawXjSNuSvjGeOCRoqul6S8+kin5UGdo2KaBQcqdvOdd/MCrMQu9KlNrRWtq/SD54L6n
QZd45jqF+lmNZMMkeKKEprqXxERSyAxcfK/7UOu3MVgmeHeJR9kN+xw1gyUa28+FaLzeGUqN6yNy
jkOoDG1jI9zwkndEf/OehBYjHnbzIXlXCLE0okkc1LtE0ScJl0IMfLve9E4tchMmZ+A54YnQ1zHc
3MUJyKnaOe7KMnJlLz5ASPlNOuG04s1hupYSYdeU1armTGWMDmN5X4rOV2kgF9AWHtfCY/Cwfne1
DgJzV+7AwZaWa8LFx+Elg5nK6VIibRIJxDjTXyk1+eM4w5oShUbnIQFxR8WNx+GJZV6kIqXW4Plj
Pg3ltQZPPSY784tTopRgo39ON1Tk1IK7+KGWgUZqK08m2MSDstwXHEo9pEfAU7cr7MoC64DfQ95M
428mtxxH3tyPFwiWmszAYKp+I2+HDc6SsOxAFbWt5vSVwHTlDCgC+ORmNccE56KMbNxAdVHcrZwI
DY0eXNX7hnZbwMTer67q2LxAz5TgClOtI2s3KH14v3y1y7zerTTQKaRuKr/stU7XrzH87rWP89Ys
7DLSn4coUn8sCKoHPHgnhtY73S2TeK7JxZHEHHNDZjB5Q87CAtOFnv2WVoNjpiaTBpgaRNrysyXs
9LfwAfJmUjtebWKU5bT1aNWtsyelp8Qe4ZpXrZOh/MJe4s1aPdgbQ+5xzQwtYyBghDx22eSsFEyX
8GQVx5NMyK0uhGfmxb7lG9k1OxeuMHlGjG4xt+8J3Ar3p39eUmSsuoLuu3Vd2pUsuVXiqNUuHo+T
mA8Z4ZvAhoVWDXPDzSCQ63jJvkdjQJvBxsiBUH1ABC+NRx1gJtqRfWBX+ZLQi2fA6Dpv+5Madh37
uCndjbbk0e/pSdeqWaaOFPhuqcu17oqJpMM5/GJhw3rD9UcKKBYeYbWS4cdeAnPgFy5w1WWMLBcb
hXa8iwIKFneYJrTvK9ikNBsmAyvlgCUBWlhpkse+rbPgCZhN61/+dwM6tIjksjdwIc1LCqYgo+t9
9ca8eLrJ4V5BKDNqCZgI42JuOGfuHzHOJvJtvWSKt5pnc4ilAyStQwbthgzRTZsjxWSQB7EGmrgm
DFRpiOzZfDs5naLZj1Erzd2U2XJOXuMiUeVElh0fkrG0BJ6KV0D++GyuQ3+bHLeQtx079XdvSf+i
eDUYlbkjd/y4+J5YO5XOIpoYRn1EQGD563PCGMEE2KqkPhvGYK7IebC5TPkjSx29ivocOrX+09xe
ujTbqWkgNFBLYhfDGEkqM9WAuFTLpf1hsUmUtRCMBd+oMcoxjoLNH5IO4/nl7GaNG82KFyC0kxj5
IEUdZrgeJ53AuwczGn2rlUG+Qz5qneteoCLNNegm4j3g/QNhCXYjceeHSlqSjiUwx2Y4Bh2oXRf2
zN0fw7RzMP6918mdjWiceHP4QWcdgm0/5Kp4KtUzdSWPf56ULl42co6jd5jY2L3JF9jZLdDrhpgg
J8Ik78wqf38eNAV27gf+k7wJ73MN0AnCYwmbab3m5m7G+hOLRNt8ZyYVm3vaPcosibo2/TQw0sks
hW/WVxk3ORhRd9UrBaimxauUEJFOrKRnSV1JY3xA/nKQtftlW+Zbn5SqZ+oiWmiVfjCP2j5Rv2NX
v3lAvO67w8UD8UuVChRuRf6lmH66fdndZ7zePXgmQ61wsCUQsLisjwkcU+957MC7sGgi3XMM1RSc
X0y79QbEFEoZgodFwuCM6cxoXgPZAYeanUB+hiFSPWGPWOhUGxzsufhdtMBQDg9z0TUVSEwzgbFt
JYuszaNCy5Z64CsyBollgKu1AbS73TYUULszqXPxgjZlM1zvxzO04PkKxyFBqOjVwJBQUxI/dbv2
F7dOWwabI50teu6ICqxG/5RtJePpIMYOcWVV0Y/2m3wzXh2aAEG0CW0kgAC4+vc3TX+Z7YvXAhmx
BdLNzPDjQpieDRcPRSeLzQGQNOU8x76eStsFF1THzPuhAEGgRyGkBTVrxG9nhoXHAt3SGBPEs/ZY
RhF9GT/jvYL8kaPIqSUU4xyqev6+zjS/D1JMCujI3rOPtXrc70ldZ7Lle1Bvd/x4JxDQLgHo/842
lNNmZF/XnaVvw3LjuI8bijAn3/Z6Y8WKqufYkmCLAbepaS3X2xkhAlXYu5IGKRpNuDJkYkxmPwsP
Wb0ItkaZQXRYiQ+1zUegRkyFa1eA65k3zFJIBFqUJBmcdtU2uJw6lmYRfwXoJUwSxFhW2qt4IL47
9H5RsVPQnV+WbKxArg5AI0N16FlkIOC/FP2lU1ufnDaQDY3lodxWnVqPrThbZO9Ne0yGN8PsIzlh
+dGtARBrurUXUi5oyzr/8eA+phNXRWWBNSugPbKLm0bEUnoDVubBGLiIwZWgkxxCVZMkaIMkP+/l
g+doVgMDsEbyZKfu4d6n0i5GG8fhKe3Qly5c3PtNg8AjyrQZe/zr32XGKutDAVwkzESmQTOX5X/S
wBqH3c1d+Izm6wCIZv075iS1c0XS/xC4wou4DWcr1tn/3UfQeeAfhBhhg6WgE7NVbUnGq3CT2Jmt
dds3DpclwrhBlh/zNljRCFqdGVYGEWelDWWz31rEOhU6n9TNMHSpU21tdbn9mLEwhXMAEQsBMjdv
qZ0iv7wMT0E+tqTK9B+maGbT9TAd/OqtpRBeh9w/ARSyZn9DE+/cUGLqTH+PDHF1FRTGsPVao9k1
A1JvjRCzj94jnTDSoda8xeQP3ZcnWp0hrCRpucuGuHOpvJK6hYKUgJnpB9MChsXfgYKM5OfxiKSU
BmKRkEq7hRb0OQZ5idbXP4IGAV4zF8S5GtLisg4OYBdtZDybFLmBYi40RgtxyNsrtDubvQohJ1OI
NYJli9rZjSOzqNO+5mNUsaPj7HMy7sjow6ofKjeCqOPB21/fcv3uvv2zGa+bqqfAzcKyz42ACyUM
Rk1+ZIxz9rzPs7QPHcizyLpfo5qfyobKondpe4XJvAV4lxVEDD5qMlo5s8y7VtEq7oP5eXwDDZr/
sVJ28WDKyO58/if9HB6nsv2KVnEHcbHp3PlGpQG/x+u4dr9hKLWXWK7ywHzR++Z8P3vGmfql97Uz
pfQAwaX0sFlclryP+5L+aoyVqLxQB98M9p5TI0xCpH2UCxIrBEqkPKQBoHeC0DKQwlA5goQD0xJ5
6bl49p96jRejObORcgkenLFVcBvLgipV+o2FTsDg5UFGNQX6ZptcKEGnLKmsyacOy2MkEf/417ap
JS1XxNdw6FSCbvGVzNQPZRSayYcFYJGV/NpMIixqr0/G6cL3BNafIj1E2ySiAayVpkYTeOr8srHz
DFR0BHXQD4Clf1W1pl/YfwvhmOV9VxLz/ttwgH0ku+VXG5uToflaF7dn0EwLH8IfgfFWhKECQW49
28L1/LVAOL9ZqS6dsBBz8SsRBwCTVywxAb3RX84C9cMC2nmr9gM+xROFgmk/vBRMOCexqaeg6wEl
IPkKaqIbMNg55arXjlMy7UzMBfsOitRcGI1+wKDiIQVhwhBeQW4/2GtqkCT9f0cLfcZ276ObxOqm
uXSUhzmlFVO3ylog3rBhi3bUw9KlyDeN8lPtdga9IYzaZatjcu4HchfePfKOquO3mudZvMtBLp1L
m3LiFnsZxhkjhfrHYBEZwS1wHXOGloCCt3CRtC9Z/50fpuZoSJOTYguS1/TEUXwkkrytz5csboqa
YT7NRU1o8Y+aweJODiYNYFYeFjBm2uW7JSr+PkXihj6AC+O24kIkHrMxRqcM4b0B5vBGZSv95ib5
5pD+/P6KLPIqFZ4VyDwjnlv6/CE2ysPgetRi2lAdktNWnUnBVbDJFFqVoZz2JXU3LCSN9pYpNNcT
piAmxFEGAU9i8rcFFZS/wRP1ufqJAmlhnsTX6+5Ci13mUYdQJemCqB9F2c9KEImTP93ytNUz3+Gm
hg3LIjngbH2rY0NE51cvZDPdg74/cd9ypnGzTilhO5yShp1okSYA4TGHwvTJHAFrf0mkpevl6F/C
I3uenm2XA9PNV5W5fh48oJ/yfPlIMHjquZADn3yixGAUjN3o/hzuJ7vgyxw+LTO9vgI5yerD/UKR
iUl1VYNDMchX07UDQhIMER6IkSvD4qoB2Xc0pluOlpGYaZiG0BXWgauDVO78KRT+30THRZLP4dCu
jl4wuRxwo8j8SQOlp1d9PMq8o0bZRVP2PsX+xyUV+R3/EAUebX+jYhwCQtXaX1NbBdEep+yodsjk
ENH1xmvTZvCBP0B18P1qldd1QGmviG05tk1oNXXoj9o47OmPPR1NBBiH0MbeGp05/oWILniHB4hU
ydTeJYfM1PTT5V5TjYLcnhyjOr5ogvjk3CqXpNeuXLhlMXRuQdlkKgaaL9Zx5dzaPDY5WRjWn1dc
zcemFvI0ZGL7HAOEn3J/9mMHVyL/VTaAZQE4vlHBDLosvJvWw+tR7u3L26Ueox/jHwPU0mExu43/
9/6Fk+/TeXNrmDd6UqeVnkvYwS2FLe9cWrAiPzu4hogMSUDK6074hEEO2hMy1krOZGDZLtE7ZmOF
x4vqdOUGBSB+ZeynfjpwasNAZAzc58oCuLnVSliRiMX07eGHwC+MLC/lhc0akanGcy0hQ2bKwVYC
bSQ7c57NJpn9jiEA8a7YmIiC1WjQxwRtGjLQP8EDUh5U1cDom98XsJFUsRhtM2RZ1ainbOElpmNY
c0OfK/0OWDgSExCUQxec6HX6fTvZzQXfEMVRCDHFCVWaiTeoBi4og6+lESaaoqkeFQNIkDINz9SI
isk22tmUQd8A5st7dHBO5fCPCNsCoDamEKpm8Hgtus9DbRYfKwvtH78ToBJ6X288n1SCoIgMM4BX
lFoFEyGxpPVeKMo2uftoY+Jrqeu8Ibk5WVg5uUBKHWDH2jZoS5IiAlEaq/f9A/bGDlwTcOrQcuwJ
6NQtki5cVi3ILRSgMqVjeSdoEhD01yalhSSiiw8DLSzFqTdV5VVxHRKBjm/O4GHksjqk1C+CXlf9
/XkklkHq5/mt4CPe4nLvrCAKELq7y4EJ2tfc9ekmqGGGq3G7LwxOboRvpUQH1gwhP9Vq4Gn8Qr+F
ryFh4069+hN7k3xyizq14Y6mJHqT++cuZoe60lUGP7PTNaneDWOonLme+ArF5hZK3+RusRpO5SAC
umR1Vluu97q8pxrfUaTX8+4Opa3iPxYVUIeEanIC+onED6NUcz7erBxPmgi8j0ZUnh38SY/f8Vrm
KcI4eK6yzyn3XPXq6HG0pyvXqdtXww4tmGcOjc6uWXwR4RV+f9QmkB42y0q/301Y0Fi5znQ6sKR9
9lTMF2LCujjEHhLhKePVHV6TkfX3FmUY7lyAsd9tRMwTGk+ZysCBx7uTvXiPHkObiWfzn3OU9Ll7
8xYwS8fhzTCD8dvS2uISK1PFy1GPbjOPBjmvIJD7RKYzSGK0t5lEigs5veLvGm69Q21uK1MRs6vZ
LD/br/WIfbXE1K19xDcrqk+paYJNin18wPMgvN0zTe3BCFq75Y24lWduxFlgFyfd5LO85cQTdOi3
gLzerg5nt8sUb8cjwPMZzKam8nNykUIxKL+5VLgij+uaNUbASJnaj1FvmQ5+IAN4B0SIKeG+gXTL
Gd+B00BuLGz0M+n/pSLLgGsD7E7jYd5fCZUiGeP74XUhdCYeZfMd/6+JAgWPQttbpbs/EBS6Tnhd
sZEzq15zQwMPF+I/I7A6ZUGwTjGbsSEmy2YMIVI53rxD/4RQt/krKzqOW3dtTbY9udEt39LWmWJx
t4KZDWRJQrL+55iUSVm2UXIlEdN2W07HDYX5SjAWlka4q0xEdC6uzvKvJIc92qBmseeZKwnfwf8w
NRAObXdU8Tl01qT8sgfxoQsYtAsnyYZjZCjFpP2jztakuZgyUv4Ohvfxb/yhjwNSs2WgJ3Fowq2o
PXDL0xX7FW9JYlf0ytKVFgdu1qV5jCBPugs61drshsyo11hMyHWOe1CEkyLUAaXV2NnL7NFwTu/3
fk+o/839zkiRYtLYCBxPeNw5Wbocf0vafm7sXExWAfZV/TsiEm3dTIcVsVQfl2VWzobPkHG29RnZ
uZzuyEc4XcO51ALt8CheUZX+mKA34lG3xYa+bUpqO8B7vG6NAPEmEFn8RTvYHgMhSHGkiIRoBSJc
Q3VxKLbQPJAUAfRW5a1WaCRB0wT2A8vC8KQcD2+CXyN3lFRO67WS73tX1NW1I/DBr2PSW0ZMz2q2
2KX2m9kXz1jU29zg16uqj9GK+dXJuQ4B39kWcyBdpWJ4H20f6xgkUrB2TxaYoxpDh1E/G0zb9nZC
+hNu8Db+9MTHVQOJ8B1/Q266wOO0fRnrbPwzD+DRirGnpGkevGjNlBO1J3PTzbIJtkU1IY+f2E9l
a85C6HsisjyvlGwpD10/PqYs21dAba6C0+8MYk64Lqp1qNez5cxKdJJ9LwY7sUFso7yd4DNPh4ac
kcHbvUODiQfRZ1xvu3L7MSd5AveuLjMZ/9Ty2om2HIr3KQKdR0nSfaUWSpvcrAPyi2FulCBysFb4
kab3wS2vr3TI807rgxhe7RBG268ZI/1Qd3ifdT4S+PQRDL+9+gdAiroE4PY2gzuSHT0RtLiaUOyz
K31Zimbc7h38nGilkXCg4Pxnba2/U5fkKUkHYUXBtFCDOyYDBI4lHEkgS2Dff+cC6ekmgS7H6/Py
akbO6N1yrR0ufR/NNAndQBgOMbWBcom/tAFw8IgtGrLwrYM0GRkdmgMO6FQmcTmKOwy4US4nOoCq
o518ek0f9JjKuoukVT6UD0QYqV3V8nzpVe+ef+oH3fAdOZLYajL4f1S9Q/eXVbQ40MdviEIwu4JR
FnJSxCQXBvbeOib9+lgmTgVZN3dfWWE6HKK3/GTl+4mONB0oKYhyCknkKahURThFF18cbFBJzEHK
LD0gczO9Uwxa410f9fkmt4A2pWKysSyMhQ2XXNTr2onPuQGZ9IDJ5wt3SoOKaalRr1tOiYxTmL3l
bsVPV5SPlXd4xs1EWp23C2TrU819P2E4PjBFFHPsRdu7TD8TdpOb7eTn/rUitPTvqSFTWlnsybD8
tNLZ47wFf6FsNrvqgOmJsO7SJxxu1+D4lrDgpkV8a1b88Gmm+2zha7jsr7PZ2uXo1Jr9czeAGI1M
fNrcES0q89aDnBmy4ZMwViWwObKvDY+uxAfBJ9lDFNfPSF+CPpYphgbPcwfdtyUSntgALe1jWbaa
/FySR/a5MEqKb6cgh7FMjtCc+Tb1poi1mgsPEylFzHL44k0JUNu1nv2D69qMOJG5FY8/9ichg6dF
SbIbk75i4duTkB9SGrtorve4TcS7GzvnXNCi4HdlvSjC6UU2y5q6JLjFcjpAVOCUQkqMgqCrZ1qS
XKrcivG/TjDyVHfvbEtuYTYJbuR0K3Go6ncMBWp2wMDYG7M1Md5bC76Lv5AsCKv1pVNLwoh8qWqT
hP9nQU2t8Xb3aEBdSzFTbKgz5mTJ34GmJFuNYHF3L5oovboqLu3xan4n/7S4T6Ft/nW1AIHVEsCl
O4mrtJgMT78duOckW/NTqhP0IXujYwXHpBE/u+ktYNatY8Yy0vr0eKz7m0W2ukKFqLJ84XLGAh4N
d2ftSHKLKNUejUjJ9hHWmy1GSro74jawsCY2jDAPntRojFe6j8S/QHjfPzF0Jtij0N+fBo70AADt
NiQ6eagw3AhvF4hAJxxJAdkFHTTgDkuGTcV1hC2XcPNzpPN+pzOFZNoclktTExq1BKSzU9QRJw9O
dUuhYmnfb0zWea3XDebro37FcLh8yuwt3uZqlSkbvmcXsQZ3gAfK2OOGwaozjXd58hFzFcRw1Xz5
1AxgPo9/47CrpcyUPNULi9Mc17RYr4hI5JzlQPM+J4qXIdcTsFF++utTm/w9OdSNFItbOe4niXuz
Rpz4+jn22Z2PYxADBnm/11q8k+Rkucu0wXTwLv/+aRwaV407fzxXsyvuYy4n24re1DECv/4vTdaH
maB/Jac7KNiBB5JyGKZoB4IdX1k4NZR7NoLTCgKQzUmtWtzulkXk61EAWhid33yVQ1ChuYe2Rn3n
MApouHBZeodVra0DUTO5Pj7QQAIHHp+3CaqbwCt3kwx2Vkw3HDCl6V2RxB7EtzrpfEkeadhtRg4p
bSymyQJyRv4aEdwGWXOCQpv4LVHtaHOoIsJbbqGo8cU81GjsG2V9/Qvt8HRa1fS5LzIMToPlHmAm
wVfEUofONWQZfMQMluEdX1ucn6S0LL5jrL0w4+h3h+WhgtzuMDqF9f8cGWeaAKZcIAADD+AgPSxf
4qZodJ5v5tKT0BMu9ZHOa4nElQna6pr24XP1/T+0EOSQrAgkFw4ePOdgCOv9TB25Kn8/bRxjgJ7c
R8CYmDyoC05ofv9Ws6YHOugsK4VYnUPMGGjVSRh6fVw9DPkCBp84V4z9JJ8Dc60C9KwGZKakeG1o
2ogvcBDRYlS+ByBoYkjoMPNBxyhYOLu4TIfNEyMM2xHL68P8wDplgaNrNtF13MdbqCTJRBGGqLcc
mDnVuhJJDOlEKsHSiAALk1NDFwrqqPOXAkVNig6bqfLG+C9Jp+3q/F4Z7/cOxGnCGQVSX5XLG0N3
W6/tUveG1MK22NLcGMW9W3hDkuu9MwNvIroeP7sAWNe+Kiw0Odh6MPbYp7rbjop62NafI437IkhD
cZ0KY92R34wSgRYehFg8aTe7wgjjcGidASX+FJc7XWflka2fyB8nhWccGxriGe+ENMdQSnYdQ85O
rInjTg00ytF5OLqlJSebvZ7eG9Zj1mUTOa31e8g5pop5gQhoYe4W+BcHWaxJZxuPRtt4W9FutTdy
J6ftkYsvSt8MYF3mf4d9nwuZg6wSyxaf2nCCbIDvIycctHAtn2kHmcts9UbAx8Z4y0j4l3qQKol9
cDtFB27bs8o+L9evZdpWI/dUMLk9I7b8dw4NZz/QpsD6EqG5z12JTlt78w4EctbRV+CrIP+3u+/K
McCu8Wbaxx1cGKUd+Ikd8XLE33wdvaoWbOLTSQPc31yBWOM5Loo2gFv3pWkegZiXL39QpL+jHKF3
HKPrgpU4oYks4q4TnybXoWBaVJOLUUZtBx6i8/7t6ZBdr+qPKROh0npD1ubDxP3McckwK7x9f2Zp
NRlwrjsqdRGR75o3BO3DdgcZ9IUI4aFlISJeSH1Ww9IaGZzDK8+cIACdJGNvncnulKRYkBygkhaM
nOZfs1osuNT8Mg+Wps3B3kr6tMQ2ggJyCPe3ViDpKMdX0vrdUwO3xS1W0dbt9xJi/9bWrjsQvLwy
O254B79WOQ6W5LWCXvy98e9TbZZyoVkeFpXoSjt4dsIsori48pqNBFpEM/7T+wyr3NhBsMhp678L
AQAKbOPZPvktzVpm/WOL7kr7GFGTyDv9QqY6myC9UcOX9ccwvHUUXIcmnk05qsJ/9gGdlMjwQkVz
You0XK1LTR/09x4O1v18OdYzCT1pP72RoEUPkbput7PWTw6KKb2wxHMil9oMRK736nObo7Ekw/Dy
TuzW8jYs8ae31t1H89BlIsBewu+VmbSSzL8IU/cbD5e46pNmgTC5JgQCa++8P6QRJenDgQpWlIl/
ueCo9Qxcgwu1hip15vUOkvyRI/+FtRREQw7RH52BJSRnvv4+IeHidfPtvZkxRZPpGb81Q1cPcyRv
x7tftaghlsKZi7aHzqlSYk5Nl5DZ/Vjh98qeBGPcG8M+cT1zU5q6cmFoemf0kjBirtI81SS2YROB
qQyJMELTPwWD2Z5i0p7y6H6KH/qJYA4DMbuihgJngkd8D8EMkVRIK7tvdGpyLUZMC871wU0SCnxn
VFwdKjcti0aHUmhchqEcHnMdQkd6RX49UmS5Yb+DBq8trH2opH4L8KRrpSl7E1BpEqcO+5p3fptb
edWCAEof7DuX4sNFCeHgk5SLA8IOqJunVo4+n3cWR9eima59SfJBUv1DzLWTodPqkS8RrpBUw/NP
v/w43srxhR3e3p65i2JiXRyKoNB/eSi9oCtQytZLz/gDJ/DBQ9GDZmDN5l2TIp3iHzNEFhVeSnap
VEoRRXVd3c52OLc2Egx69xIw18PjR/RjXs5btJPDoV8xylVdSHYvLhVpV/ohtmI8KcMtpmd2ljTq
YqSLfr5CDEtkvvWlgXIdi1S6XZIBdcIm2EcNLIqYDfzWIrsTtbcdcNqt2HTNbMk5Cj4z8CWGlNGD
TdtFvWDwo50skUzDkE6r5DmYQ9UKohlwIMrhvDbTimNpfcOB+3TQEdSGn3LCNsxYcVGxa3gpvv85
YM4hnzdbwqFYGLjH6dZASoL4+pPPB72gKEBsaCXWAvRN61I3Q2EfulSgnp7vm2sNfprDV8WrsBxF
X0wVo4DQfgcKWabJzSdci4iHwS0CXMZHLZluSsC04/a2whRMcV9d6oG+Cc9YHRcK9GqUfI1r88/v
iybx153I8rqqL5Is1oRZDBh6HnH7kw7IZhOqKsWmWbiobA9zSa0HNWnCXfylFMmTy1WKN58Nia3K
bQvpFmJbXCqFUw70vyjpdjSrmwx/YB7OjQpD9ddPgylXhV59lNR8XmP4WjCRGnIFXxY5cPA/SlTS
7OveDVFywDKiegI+zlhIcWZkYUgHQOVxyP3P6N00chtrNIJVNRK07W4qO+F/T0S/4gb6XilSKr03
S/jSLER3xUc5c2tEe0+LzKLe61my6pbk9CAQh73F/UUFa5fkP/Fz+yVQRp0oK2AQRpheY9dddp9Z
2bkzCm7OxmSgjuaVl+R4JjccRpTPhHK/IzukqQVHJAvadtB92uLHzvOHaS7k2AYZWZeanvcLAmW9
+bBp1GE+IdUX39UAoM+hAOPKTpbNpMtgxbpZYWwg+QuAjGrXWQlmhbdMKxBbtY4OB6wL+CQ63MAe
uJH9dhSSwsArPLze9Ze8D50AOUQL+dQQe9B4J1HLioGGkf/SLGsr1kIVan0TEDwHZl7bOo/Z1Dqg
meUienQneRD+Asgd2r7mjmvheCbXJrWDFiXF1arzp+eCv3pVlNRh3A8q3tYoKXXHqEEUzEoRoOL7
UEIy8qYXEBXh9v/QO8z12CtO2M6bD+hWWUQ+l1Av8SVsYoLjNBX2uyUERUWmtAaYix//ABkt7KF4
NjM4Lr/XYDJk7mg7e0OOxxr/eOWLZXZQ1SBYzkbNJQrglbo4wJSB0qFgg4zPd7YXwJP9TY8NnAzM
MijJpZ7Bxr5gXRtlShU55IiQbVBT7U9GBvzD1Td78AIuVDt0SeRWnRf5gbBJ+oztW75pKzamGCfw
ow9o4OQgOvCStAgfhetPRFc1xGjSV7MRE7yMxMbmI2+H4ItAUUaWnQtHDOa6aF/V4+owAK9CnoQk
jNq1s8kU4OfCsqOUyF/HzoPpigZUK1k+D+GRwQlIRTPhfrS2OlB8EL6gKyV0Zqt6wNPyetojKAsL
hgbcKt5NC+Zvlf5HqeAazMm1YSm6KOY+58td1EiTPAMtdo2GBTmt/69kCqC7mhWfpTydEw+7Yjx7
mTZd/T015RWMwkb4mTxn9rUJRLwWr7QgXgQs66lg14+ygVmlyPEDJR0qk3tmYWu39cUnrJtuQyBY
pgMaevuDzyfv9i/yQHOt988b9PA4d+BWnWOCHs8Q52NgYdFALRlW+qRJTbIVMRlShJY4VEDVxHG/
83CLeFGT0XlH7UuLERaG1G8zSULTTDGCFX6IgDHkA5dfbVMsvjPPT4fNsDoTs5KbN2uhij13a0Ai
0W/1oCB6ualg+NTsLqO0IlwNVFXA8hLLWbjJTehnOxWdMSNB/npnHCK/4KevBPRZnv2ge08fdGN/
nM68a0ysTtazubgdKfjnphS4AhGsE8/aSLShN7bhl+bISugiqCTF0WIzMePJQxpy9u1cCF4/zMGs
48vlCvIVmye2iDuFQP37Pb0dr+94SRKpMir5qQ6ZkkQy2z8rjtCNt0crLlykPUxIjfkA1/BUZomi
NsyIlvd+Rf26h8luiBenFpxs6ord9UpJ7Rwo3Dw7hTCAYLl4ErVpWr/T3QjUFByT/+4y9PWhmwFe
E/nr4Ftiq0hAWb3E4T45SMPeUn/3r3Co7um/U6WfH6TO7dVzBMZt7e9cY+A38V9vyeGnbsE3P//p
EqcSmhgpfhaAV6X2Gb3mD30AatFi10AxfqbNeCmI4KhAH3T0n1tqqOYAcmCUsWaTQGEDiGQkaLEs
dZNCA60sH3ZNuHLHNpSFe8xm/0NMUxEuew8OYkbQterTUMJSDuzCBqG+XK54gWsLZ0RQccKHhMoI
k6DuS3kp+q6OIZr3IZvSAZ8p9lpY0WeezXbZ5J3OafoCzsHAFi2WETNwnoJ4+FChWqCteCYYXWBO
//bUvzEDkd0kQCpBu33Bk5hR1SgucsSA6x/aFqFwY20n3cnNrpJ23hj018Z6OGh4ptsk1a/p5ZpI
RWxzJvcc4RZ1n2sXOXjYzbDW0cGP986qEs+1R2jClEXkJfkGwXFFs8yrJ4f4LGyc0TVTIIm5Hm5s
eYwvIbEl76Lt3ZZXLpo3AgGvFFYovOjY9j2LrVJn7/CGVaBalncJKbuFlwxIRXgCXLbGEIUtvZtE
kVPJLttNQ9PH57rGAmn/z/cOrqFYr7O70FMO+dgZCfzL9mU4l5JlK8WCKRgivk/vc6DPrZYY3n8J
KV3RSS6rC9KHyhgUyzuSu4j4zP67/jWhdBCsSmxQ3VGCDnC4G3fWJNi13LXFW0qb7NL6EH/WU9dA
a1Zz7NAaSfmO194n2qoEpjsfLJORWEAoRe7rJMOGa+NdbyivjAg9muc+g54CNhB9blVBYaZOMc0w
YR4wUTwcdwxqGTrYI0y2O+WoBOyh3S5jKG16HDwWgGRwUjcGI0eur8QoX8p3tdihRgdw1754ozCG
tnA05qqBVZjgYqfw+Pz3l6KflfCqkL14b4RbxlIEXGN1tHtWuF3d6SvZnr0yF1phgv09hGrDvlrW
2a6Xr4f/zMI+OLzwU28y9mL9U0+bMVNI6/XQk4471/2J/J6OXagnxQ9QJgXrs2oGycSZnQadds4y
a7kZHZ0s3Q2fnnj/2efOVpnCHg6eVhMl1wW+Ov099Nm5BXiF9QkSDvhiLkqSrnrG1iCnZ2MUtosH
d56XflSlG7X1xH0LVwTVxrjvCED1A5SkrnG+VrUIDeWv57o3NrqelcNZPCK6JykuslI61xuc28FI
m02POIcD4YdaEDyo06RcqKI9L2pAdKR3rnQloZ4UFdonVQNGSwUNl+uKEty7AhPXLljwmKW4hvoH
nWXTsiFWYb/yHCMXbd8erk/kAvihauV5tr3gVUZOw/cqX4A2/C9Jqospv3U68VRcCJHEUbj8Rvtq
vPmwR5f0wOQJveX3f37667B+Q581jmbhBm4QS3lYKlW/r4XRe1gUhcbKGs9eeChoNFCfhLKLY8IQ
SFIuH5dL8sfd3ZYw4Mndhj+H3icvIGwy7FartyKGTP5mOt0SODIxnu7TzjC3I3C1fOF4yrTQL6TR
+27nFtWOaF0UCR2317cmUMan8n+K8nsnTwUUxn81hdO2U6l6uqSCXF5zJIkO4nq0LAxFJNu1Cnmt
sZS5PAvyyP+Ewkdo6PvsPSsgpdFPvC9pzKK1VUJuJltfz41TbLshrT9WZxZcQdnNUmGm7CDh0KXK
k/hSiNEdTqFIeAf2B4codmNqTO21jhYGf2ONrGPu8qPd4/mxLAp+JYAHcRIXR5gSOVNPDpfLHWnb
MVnqUofrdyf+DqNvcQgJNSM25ucMt//KULXpo8L1KhXpLnzlrpQ8gfD3jMDXTzt3Yvtzp2bF6iBK
ASTCW2xCZQp7Xr+wcv3Fc8mTWqggA7RYjnIQg8SxEk24QGrH2AH5yQz1P4SzKXjTqElgjIfrGx5g
WLwoGXUC1cahGkeO27LG5kpfQHCrFzCoZWaZw389rZKqOGSecSc/9ujxyutjymU1zpNfQZjyz2Ll
aj22/UbiSRaUQtlyM9mPX4A0e7qImcgQK2CCkUcfJ6dXvz9eG8BPXOGSUSPxoOnKcHctPtjb8OV+
RnxF4vlvJAv3oadrkCspuWpEvoFsKyRarlt1qH5wGoHu64aVTiwFof5RcA1ae6BmNVa2swmzkyM3
rp7kl4PgTwh1F34M3HGldLf7MqC4C67q3Be7v5Z2Di/rZ3AM9xSv5rphCrP1IaJmLhojXfV9i7BC
2dBH+EKx6hsi2RQEZx9jt2tyRVJ6ZTP2j3mEI5sAk92baEvPyOa0G8H1AN4U8I/RYO49jCcOEH8y
tHgxb2k6XBiOxn+/g8Y/VVic89C39b5fXBj44uf+4KmfVE0tzcua1ysO3ylO+zbe4nACx96qbiT3
1g7dFzhxkRDbxzA2aqosa2D577Wc6NW0KhagLPiuUXbupymT0JUlOs76pW7l5QqUwaImQgHOoXhD
gogJkvDlf8Fedjk33TIEA5tz6gruCTnf2x/cwF9AzdPb7Thv96qwZDd7NnJw93+I1XuGT1c4zxVb
Fgu9FoQRU9hcgWA56CElJCer23TiBP0FKE0CzdAI5ECpM9wFA8qrZb+K7LYep8UEZUD10XMmnAap
cNe63JrRB6Q6C5ACVq+OaVM+zZwnpDBRTOKV0GQ0kVmqF+MH1+GhKqFChJSLwvPlbe50OZztFcU6
gCj0YUN2ZCMod5joD2uNEHU4IDp28LHp11UZ9DrIMtK+ftgeXFxNHLIpbWUjr3/j/UJK/LAVDrWk
qAbwe9u6tSTR+fneti9rWN8PfQ6e5lyNneCW8MFz087SIvxKJuPwmUMp8VvVTElzPWClWEabfFPC
K4vWbHi+GElh9irX0/RZLn6+svFwW2I73tWa65h3PMksVqbHPvZ3W1oIfEiZXxmoN0eNulv6wz/H
C1VOwQdVytU85fYE+gm1mzOmfThwF00UaxNFQ9amStRK9n/4P+hoIgt9wIUE4lhDC+Vsl39TlFT1
kJfjHUA4xvr5xdxN3aHUPzgcvbZQoDJrDyMoWNbHwU+xMtnona3pfZr3AyUwvdRx907OzP5dsE0W
tH2Rb9w+uPRsAUlT7GQ8SVFhiJygMaxeATCsbKv2yU4e6yH2TwyvUuz+rMC6sjdbzrZRBQMOx3wT
LJRO5lfqqVvWryyebmGrqbSsCTD7CL3DnEOvuxq5reJRopflTLISAWm3X+2dgdRhbYXzY+oTbVLD
cA4maIn7AuDMMbveATXZZf537kU6nNM/s/DlxfkDri1JV0XrUk0dqLZ2ILt2eonlO558BZurlbLF
4OQqElpm/VnK5xoOGc1NqBd1p9H2xFWBwa4Y/ckM84jZC9fEpIRAW/I1W3klTV+jTMuBKj/JVo7k
u5tLTpmVuMXy4tiSJHBbp6hlFoxaewM4AZc+Om6ZeZuy2N/BggpNkVriUYVpxWsifWECyxKIiKnS
BfIhK4Tud0MDKAy+UpsZYdpCQfV1lm/g4XBH8kfFvxSFZS807JLOjDRRcEpmFHyVvKQTKovdQ8yc
XLLOI5PkjNbXfsCPrI4oPWRe4rZOkQPLZdKhrzQkxke7R/IiNt8DnoLp4WB2x5/MpOp4w0o1O+7V
kjTbQiG03vTWOSGfyqAEFCiaJCa2AoaOJyDiI3dXaOgCdLHNWJnZSp1rBLXELiubFVh1oBRI0UU8
kf7Al3Pg8aVIyAxEN30i27oJvy+lv/UCR3F5fu5R7qTdc/5iQ5Jz/ewLHd6d80FKJ06cdrkoEQk/
d/i6fZaKfv36/DttmbZhqjqsMrdXqJi13AeLwg2gTjv/n7PJ0sXTQvwd6zm/saJ0KiutImCn6IWj
VFA+dHVI0OYlkJr8hOY8ZEmf50NoVxiT9kbSAzvKAPvDDsDA6yPBtHnCQ2eY7TMwSKk8sYYVB0I7
9Sk1iqYV8qA0rn8mxcsKcfoyq5Nnqi/bzP+W71+qx26vzcAK/ykgPRj5IGJpNikxs2foG9rO+2B6
GoL5mAqzgg7/1xo2E9+342W/o6ytvO+FkzU6EnGsWxlqZsPnu+opanIAcDzETbDUkyscohXVxaxh
eqo8So1te2dO2iA5H88KGNuq/Ty7J5BukFXuFMbird8iuCadXS4zA4p+8IZCzEB5SeAnbUoLAcCU
tfsPaMiOdwnjN+HdC6x8hQYWDAnuXUSUazdogyjoi1L5lx1j02GBIXdATRAStJCWZh6XJnuzY0X6
jLl6qgoNmyMauiUNWUdBMt/EDIuya04SBrhsz+pPfxScw9fIFx0FZwlnRy06VlWFzHmI5SIxh+Fp
1fR7t0fB947S+8Bl48BCkTq+7+8B9orKJhHv/g8RdMDBhZjIxtDuieEH07zYlYVD1Iv1RI0osPEq
4z2/JtKazfJyvnyjFsJMhV5TTNniIrvjdPCL7+FsxAy/XhQBA0RZDghP7257hXDSrkgJSbHOZmt5
nNYRTjRJHZqQSsLe5nyhAbCFQap1WQ0sKKbpXC5sCstDxjJBpuwiJLAPxMtokJ30RRZn+eff0TXt
GNHK5L2cnEK+VdhZfL+VwVDW0iOF6syIQTuq8HPp+DMo9e4ECrX7VhN9yFuhyxyc5DAPHfIOgNKy
nfSDWXBUKDbwHs0ekV+IH0kvNXpRzlo9GcbAhea1sMPfvrsjuwXRjGE4BuCfDIDWFsronOYbOE6N
V1iSsjA8hHJjHt6Q/4QrMcit1dcK63PcBRmgGPyMWR2yDl2djbL0TwoBQwfRIplTIdubRjKRSlQa
ARomRQwyjZ5ODL/71B8cTpi/Msq13KQ66a6sw0zQADCZBVbb739CvnA6wIPRLwdu4U9DBBX92biV
Vb8wEZeWwB60JIjc7jPRhgWsI4EsqC8a6bvqvyJHTpkg28mIzrhG8aS/gbdwpQ4KhXLF1svRIpFp
Kpkp/ZMOc/3r+YIQIngViLcX7a5ZbVyO4+s/eMtQXmkWtfpGRc90IYlbEXEYXbk/zpeQvOhIHB5g
+1fApWnOtWIBaiAUA01cY22uUkXdSWfVmYthNNWewNPxMr4VuJp+Kc4FxhAlebfi48sIBlIYbvWy
DNdmu+R71ompmTgu0CeoXOz+7w1CJa68Gw2quXNieCpqihWDBi5edGRb+YNtOhDawiFdFXyCTsdo
jITFFfQRsJo4Uyv/lUdPhMRC4mB2R1+0Od5o6uy7+iIp4lOlwqkMUTyai0mH4G9ib75NETC/nUP5
j38U0tGhKavlJ+BOtlgSwoYrjJ88whoE6SBBBYlimPJGldJ1hHY+iuVTTY6ht5BBaE8ulUgj1IfO
TQc6xVfc4lm+QkX5ozROAkGson8NyaxH10KYTU+K+M10aIZPs82HyiJ8XIULkqOkKkE4vJxbQmx+
yAbWHWPrQNgHR7mP2nVn5JdD5CItLMeznaJFmPi4GdLEzKGhBjbHRj8Pkhuv7FjAnnt8RYbUSGOf
3V6pJ6JWU4g4O4qooJhX1Rozw30D9qhnvymnV8fZtvMpF9pY4NRKVvFgjmSSwBewhnm8qn/QiO/Z
H9/y4lVSnfTj2rJVtjhkxJCgzFNt0yY82/ZbCYN7vsZGapxHdyD1v+fzuJ85fil8Xpqv51KPaul6
FbNEHr5nfIOOv5j1YsVPrPxAv9RLMksGjaDD/4CsBVsGmrP4aKzjmh3MA1GMrx8zUMCPTix2WMtM
PjwIA+AS38guiga68c1udh+tNo65WpNRZk8Pc/sqd+fl8hvIr2L9mY8+yWKpefnnxwShpeHEFpUH
QU9IMq4iqatRaMNEWDzi74c+ZXUkF8eeQgDlEV6DKS7+Cz7BkF6OTuGsnyx7kowJLDL0MGftQXL1
sbssOWNNZD3rWPlQ3ERA3lbISFwoZtrjgamyyBnEHys3gXPTVB09x67A1V4BIub+614ZsR5fZhBy
GWmmRmIfUGFfHC+DV/SK7e6HZrmC1LXoI97O0fHUDXLIw8IB7oYxGaLGx+ZnIpLWF7QyqnLjb5Xq
4rDNU0EiRwysZwx+hLqE+Ud0ievrxUAQuLoWPjjlELB95FJHanxruPhdm9d6te2qjn6u7baT786q
LhleLyAkSvMLQPFkXi5TKE1rqE+xXzKgvck+7acAQuDAn97FvdCB18P27skjaeC1luA5Lko5jDM1
wZYumP53ibnbKmhus91xfvinGzk6PVZOmx5gHt5JO9wYss5ISSGBlSp/6C1WAxgGS1WsvYMJZs1d
PDieIAuqegHJ/jkl4LOxItB7jUYavh4GN2jTD3YHxNqCTXlef2jCB9zdM+mCpAXA5I+8h907JKwx
XhhoAjJNw+p15JomUUbiwOkNjtF68b0P1T4bZ4pSScbPohO6Zff+gatxb6wZJ7xQHZCmcvnlZiFt
oDokdfLEqJkQadd0kJcfxS2mdrEkyVSaM4X5klkVxSGmQTANyyBpEcK9OO+oeLbtMzgcocHebfQF
pE+hR9Uwrnq/JPYQR/VV81QugHEEGRMcfZkFqNiJtJ4g562HP2eIpaNeQI1eigD7qbn2El42H/Ne
M8LWwgohycohHQa1XEZhmwGdeK9QpiifVrOfNUhQM+fMxH4jr9kijlZeTXMUl5XLjnNjeRUbjGVH
O7k7Dsr9AsvtdtTyVy5Amd87sVZ44R+Zaoa7Z1zDeY8T1ek2tYzoxokhrMwms6MF86HifepNzWRw
JBWOaYp1ImQvWQ457KFr/6YqGYHCulH1hTVyV10rFOFuMNSC4RsPf+sKKKEXlkh7V1W6fqOY9iyR
m8uvlab7sC6WhFWlUq8fW4rEZH2NznsHXKv21WclhcrutjZsEct3aGrE0/kplS6QQZJPB9PGZKst
tW2SVdxP+nBFtV2P1Zk+XGcHabBGh6gYPe8QV2EauN3PygxKWdkPoNgMIHcLJjuvTurin2WEurQA
Zhfp9lXCFLJy+eH0U/fA00E7ajfPvE5U8nXNXj1guSRuVLvLYbEXd9Txf3bfIrsNuocbk8mUQcJu
N5JOVAF3/le26iLjzUNJ925MTDcznvH7Qd3jbyH3hOwjwlenXz5SJ+62yJ4/mP5S11Ax87w447UO
Ybex3sF55+FQshkSCApEA/7TfUN3fYMej+oIVSldpeT0cbKdmFoYq8rzxYo5WVZlaytYSAfmmYQ5
qsa2FK4JnfL0KFkTDKaT0mDfFOYwA+TILdsKR4e3QrfbAEjkPgee3U03dpfdZ8sTMzdC8GY/wAI+
aFevxlI8MKPq62TKK9Ig2/f5uo5jXhIdP8Eivd+Zr8He4jHaHm5Z6vC4WlgeM+giBv6ciQAsjqi1
ziyRvvblTGW3wdmmRRQYa3DGud2RnXKaeKLizMLiBFMoH21EufkrixXeyZpBGnLncByafcISDC/5
FVEShGAaza2n9DATRYsmrr8kxmk40ZbROgOtOe0PVwvz5UyBNnF6HEcWLWCSSQdNlRB4XDAA40pN
2CO2zxJiIHxR/gp5pKCLN01Q2ofcLFbMhiMaN0RznYr2m4c1BKTbsBl6y1A6AsBfJ8vMgTzajvTJ
V3rRGkhfsGGWAiCpabnB1je/cjw3zMmbFafLBQ9lgioy9BMFfiQnQF/vx21o/IwRUTjThVYMb/Fv
6eQRDkAw+ItIMzjSTXDyVRz6JoO/OvKCKC6pSopJuRNkl2Vvs7xaJtbEgOEbVeG8KLEHZlokkxRl
Wwp92k7JqYaFiVb8EYYrGVQNt2TkvPwAhJD+UOkf0QScwWu/SgAlV7Jx6vS5UN5nSmpp8xtEvJGX
uUtBKMPSf/mGEnJ2Fs9UI/yZ3sNObemOzMwUZNRUk6MFIVrqfU5W+wF1b6PY+rQBKF1sIHE+PEJS
Wt6SWw+Weqvd963DoS483mrNMbbrXRvRJPFZMfFKdej+rKcBIqL9ETxYDkg68NGWTWoj1WOPgKI6
yqxiPPrkb0FLh9iHTj86zz+BPg7K2Z3OcmaEdTGbB/WAvC6lx6TPTQX7ySmwo8R80VeJzcfPoHe3
DxVEsYCJsso8Z4U8o/zj5io0rtY0VfEGRT0P4iFTRPVWCYJO0S3yMItoN19Q3U4EbDlZwYE7r2qP
syaLEzNIzSKysoS73RwbhMzJ2T2im4u/CY4MMzlv7VhInIEZu2yG9a9K4kkm4ebIFU25QLAve/1l
zdpan6tk5ZQQgsA3Usbrs+NAWXZUvht8WVbL7gthGfp1lteF39wiyiXMb29cAV6z6XdiqMyTYO4F
YwpquEJ6V0W173Pl9tNr5EBHW/oOKRdRew0DvMfG9ibwrQf8dmVa3mezEDupf53YCDeN8y+i8MV9
MY5VC4HAiIt1knMpW35v7PcieLRFcrck0ouD6WuJSYxCZD+NFp6K3SyBUZwyDCgcr8I1AMV61eLQ
Pk90d9vZcVZ4SZH/qH+CLawD4FUn8HdmTluHW9tzGZCGbLXjhckOVu4KBbsBqQwwXAEVVYfnOU2U
3sGoS61+frrLgAp+d6+clw/9ZcMaXDKu34JdhjqZIhKclnPSyCsawp0rOAwiv5MTDTpLCShCGgEz
7zYulmzaClb2Ur8hguOD7ystZvJihXwTwOp/sAxcGMx3iyDohe/r+TsIAKABX9cvfKvgHg0L4ZCw
Cj+07zj1UYJfOesoJjo0vUU7yBVOXX67Vn7Dcg6/qmNB1YnobGuOif3JvYQSAgBd94VFTDUEmBCE
bfDcXItqlT3D9k8384wsJ1BeWwkZTZTK/as9HohriCLN3Gdg0ebXnKXLGg4vbliGUbnw1joM91wW
Lkd9/riosi8S4qLCVwfL2nK/Yq3XR/b14X7ytFn5xE8d+H3YcW7Wasq2wZRrUbN/F7l93K4fscQq
KoR/dTaOKFG6Fn67N7vjQ2DH2KvodCJwK6bbGHO7yalWIxzXN9CyhlKgOaRBRKhR2gIGgCzp9PjD
DcIzXSXPNBVH6qpJ7dm6xz8lxo/KntZhe7DdxU3kkJ+JWLMMpT7V08+/3HOAvw4R4AeyA/9e1bgZ
mBIqbVI/ljumMvjNhAC6Vp/AFrVKF1KUDnBjyb1RRSAzEvLQh5F6NPEYQwB93iRKG+Il/doVpL5T
mT2wSoiTY/3C9SQ8FM6hiPhNLByDZmj8roIpKnyOCVwlOzyZ6KvAC56DiTGzmrL8O/aNShIHUXGa
E4JmiIh1gz6S6DiRxyP2jI0vjs1apJp27SNf++RThaChgVNAbNdmVMEgcptoreATm6fMN9gG3X+E
HElXVgUFmtWdtxm2vLAeIhoade7z5+6H4rp2hIcHjlzKcCtF9SYcqP/NUFGQat76/aWg6IRG4baW
xJOeFqxJ1/Z3LyCPknf8InPCNQkLUryYbgNVSjoghyICXULMXa6lRiyVjfkOGlY+5l9V1goFj5hX
R8W4SFbli9xtEd49zpwi0HuzBfM0oOxA3y2hPzVbd78aqzw7NlNH8qNGmCJYquSkODgI6XFqF3GD
Dytp5+NBTB8dkVS7VaPdg4iHgV11hz76a7J6lhQuGgAT1K3QtowKP7BejP8rR4yKUlZGOdv4523z
FiaeE5FlekFHWDOoT9Gum06C/WXwsW2rY2A8gRHTQAvG5RQ2INwzTwbxzKTxeVdTzfxs147o1/xF
CcQnD1pqtcMNTi+SMcOJS39ouZ0gOn/9My1vjjNJcT8gxfEp3saDLseVtyTFXIfC07tSzkM7sTY1
Nuh3IneQdYNpHxKtsrZxG4QbkD9hteWRQVmOYeapZMOjjjgGXvL12vrhoM9BVbzlypj6xXqgnKc7
HCWg9ZN6ZTMf9CISek4YlBCg9FjSEX5XKIXNKfd+M6RNmTa9XnfeOfRXaaST962bSe0JvkgaQ9QD
Edun4mVoM37Cc8f52yo8qgUleOcHjd8OVXuwaSs/EH1Bq7z0ODEDHuJyx0r2VIkP5Fq1MYUpHSxS
Z9ksLO4v4nvWA0VtQyrrcrR5Z6jSssNMjFRWGe/UOOUWPiozCEIokSkrKd523+S+ivDCPfECLeNz
aMQl1wmIoPxVLjIZbnm3I/EoPGo+D2tSXzntrJFX9W2IgrYsemsYdZnrYqYO6uVYLOHoMbKC7o7x
Ra9j1m9wLY+WMqlLbIFlCAGiRQVSvYa7QYRBsCKPi7C0KUcJGZ0hb/dfnlv8wFi2llOsM4KtPxkJ
9Fly3aGmfeqY6fSIm3eI0Zzro/nPtClbEufW3NLW5mmrT7Ia61q6oDIye77X6Misbb7RHlHZXRJa
Djkd3pZx2r9EB5Takd4N2SyJO6Lc9XdrnUF4Ai5hJsf4cWSYs7BPKKYBzlOWtx5Phgk5Zg0h+H85
Yel+jisKSXvyiNcVx0gxOEYDmcOJIuH3nd0qcla2qbj8TMaeqXW2eHfAyt6+M/ihSbtngYQM/RB3
aMvR1yO2jqaUKgYzsmmOd9FKMTp8jwidvA1woioVb4phQllPGf/aGhWyDN1vQqT4SMalUeskkp6L
AHpQoq0fvaKntyyI+G4unEmYknFjCZxrXIvuogbah1j5xQwmEoHBOFvk7hFXj3xrTnH2IrakWd8M
w90dB3aIti8+WPyGAFqqT6o/pkhoqJsVIVv5RnsH5wb9V4o1xdXTRc6mrGzfli/E6v4DmTlif0Su
vTzjgUcREluZEAZmqso9vFPQD0mtBer0iIyM3zuYryLBvruBW5P601eWEnnGeThhVxbu4kwIcyMT
7MHCLYmbLyQ6DcNQ0L1Yyk4il2ilxRwT3S8QFEPbKDR3K+P7eofcOf0V3Hl1htKueVF/ufsUDp1d
+QDA/KR1Mm64WpSrUAf/RpekXLS9r/MCUJxTohthcxdg+Cc5+5rn5889iGrVk/+7UIOMB+Wo9wt7
9xWyxy1gtdbBdQItESww2myAbTUX2WZmmI0T7XbpFe+tFdGnkUZEHkDvcMpCLV4e39f2T1/+WaAY
HqXL9mmzfHaXmQ/NqI9ZkQARTR0Rj2TV39yoNoHga55PQJNRlkE3hUtMaVVqB6OVRbY+yhAI7KHS
rvMsCekgWj2cbxqqvt8bb7NX9fmziq3pWlOdqKAafRcN2jPS+LXW97nDFX+74R59kCzIPkEQNEzJ
DlJfUgjlJe8mZ9HeCSXlwsFKrpMfGGajwcXKwLUHrAi3VxlH6HYY1uglDvEGe9mb3t+uYu8uMxuj
JhDzfdzZdWyDu/NdJcaQ+IDarHRukT7dgZzDxBA3Clnc80VldLB0qRhwJaNQfAU0ymXFYQ3DaPj7
D7YKeQyyzTSlGYyEQ/z0aH/6qK4c5KPsUeB4QbCNWcuwxl7t8hYGaqt07RPcsq84KPCU/ARphGmk
1Ym6hWNieV3EaJi3JCJP2FKthg6JyO2z3lKbYeoHM8YoIzDQ5RHy75+k/EvVwkr6kGbfhipm5wCh
eqe+a6B3+Fv5xlruiAL/6XaESSqWq/acAefcCxsO5urTsEVect4qw8vCYh0jFn6fjTNdNiA4evVv
fI66eXd3izOnmipRnOTphLa3W+FqssltSi94GqGO4VP8ToDlWTcWOqHzBEYGAe4nK/oOpGcDrpoJ
QAF8CAN1GA19ZemtLcNa5mHsEqrpHJTHsjcHyxYzi8iFTZh7qgTZ5F+mJCcqOJdAPPyAOpogr/OO
BwiKlKoIkGr+9k6H6VvzBYCVlkU+uhwdJPcE7gAJEjOsfXyopCouQsZPiQVLulsae9hddiNdPHvo
MuDvyHosEaR/0DxJbYyu3YGkRzeSQozDbixQWwQiQ3WfJYswHU/kzTafZVo4mFxID6CiP0dJUFPN
/6U+ViCVc7/gd6NtJC32vJBq/TOrKvP3DrtWKnSwt6ft6J/aoDysU6LyRHoT79mkWqEwcflLmeL6
M9RrslvFslZ9l5rSxyJ1N2ztS18xAtIfw8t4lmsQ9LcSMV5SeNtm0KK4mE5+PM9e22HKI0cRATwr
bjDZt5375Mm1o99gR8PgRl9RgZlGc/8ae7K9P35wJcxdIxsXQRhwpQdBFISRfU30xSNF48k/Bf2f
/CMUxIUuPbgcX/YqIxpu+SBovqu/7AZnUUfQ1n9L8zrZVPRozXKgjkCfRwoT49mw6B/ws3GW1dWO
3kb/JKv3vRjMHFWI4t0ekQm9SsOOPdRerVB+hIYTSOUh8K6WUxQDX+kRadibQTm1mYr2j018C0zZ
sjN9EsLHG+8Hki2If1MRCkBd5ZAOLyI7fWwLr3hhal7UXi+Qlkpyuu5Nzx8Zv/w3rZaHCPjr7anx
xVBnuX5lwWt0lfqMIjrZ2IpAsbZYPNkWERd8lelsjS59GSutOaJdnn4CG+RCjR5sSESUPXcx6tDD
bDITva46Ap73+VUdmRL1H8Hwk0GVzsPTvm8nWytzHsyHk3tWAPzUhjUDzWxylfUVXISsLtpNJsTA
uLH4IQF/KmeKK3QcI/+12FRLjx3ce/NjEiHjxyDsgevACJDvLkfqByMVVERmD7LUpGVopx7YqksB
U8kpNOJxvwEeDdCWZoIhgIRG/yu3QKo12pZeQtiBx+ccEe0+7lYeVGdgdgWs+s5JvewK7YvlL5E+
VkPkVWfbRsVtNSoHDSfacZZpiYL0HLxqyFB2ftNVwY7kyQyzY/0TBUA9lVOP0hOIAgpjO1H+FvSE
XI1Xh8ebabtC87MQSpjjUMd1C363QGMZIVEoJzMQJT9NzZZFAqCxtyunYLYBDhqyhCnLg03PU4Hr
wS1coJiiSw1xazuSa5lfhyF+dn45Pcr1iHFziicvFOFz2gnrIKVxWRbfU1NPaKWzMJGDUvvRc+JO
7zZVytagrPsSVd13J6S/+JASjsZnmIryjmKpIkNBCJ0j3kBjj4axHuiqdy5coRf8OQOOLCAJ3UDb
t6SKyAyoqYRv/qlVjSm4Bgccp9KsWjMhMZBTTPk9qKuBK/VY3rUj9ZNWIqBm0VTeDyUNalH5thT4
WgNKd+NP27h9a1jLTg0McuWtRbZMa0X+Z9LTrT2BSANkgEQP4xgM6kSUhYwTC0/rsfaa5TrrOuaP
aRfwTKcuTAOiB+3XvYj2uOEyODgKYLdEKCRbMzYhlSU29vD1V6uTtP2BGjco91eIaWQZgvKw4NgD
q6SsgZWMJSUbfv8K8NaCYdPFgxaiH96mqRjSmB1lMTengbEGU8RA44uNCnRR9OSIWb32p3CUDeR2
5C8GuMtw3plriUeka50qmWJd8yutZ/zEaI/uUZzB6BUgMPmhwA4/+6LBCV0x8kDShD5FiFr8IX2v
0dCM79fKzPJ7lwzwQxkn41fgphro6S+VBKqriPmskQxFlydeuOY6WNRLW9mMtppxjVU6E701Bh5A
6Iig5wFiNXiAIeqIMLR4mzXaTJvre+Bf2hNkDuvVPWrvrKmy0f095hpTbFqAyMz10GYW2tiGE66d
BlMxKz4SEZoK4Yw9slRcNpMbV0fNPPHYTbQntcfoMgm8L/BSPbK43GEFrsNoIJDtECeGu8W/feFh
CVTa6Y1YIvmoopJZuRC3eo8zTUAQQrb/5H+rvfz1BlCsg26XlmI6t72QTR8kl38vhmPywmwxVB9d
d25CWPX9Uzz07FeM2qrSPU5M0sdJtIvylDwUJPM3rggAbIw1ceJ0cuE947qdh8vQNLchKjbHF0X8
cgVV+VBihgd83mCt1BimUbeykzBt+BIkxqW/VtwqNAPtH82Bc2xNc3xOwrZJd9CYFQYbVjDDoFZs
zYam13YpVZQ5AcQJ/LP75i9TLkZ2BVsgxOJ1yBu5if/8d/sLg+7+eDIaOl3gACarizvZCgCqKb2e
uBIsg8h2ZH0fItJjwJC5s1s9U+WgP0B59k7GmLiU8OHh4sAw559luDg5eu6BOHnstNyRDLSxi0+Z
2guu+A6K9IzLsDvzj0L7T/JE3Ju/ZqDnyIgSkTrzqhoSTTj+5fg1je5bj2Qa52nPjxR2vld9NTP5
qC/JhCHxI20kZxVtiArhWwq+WH4aZ+7KO/1wOTh5kfOteUmCBzO0MAlAU4sMl43Nx7xfeQTJtu1i
KGuV+1JLrtGaw0tabHIp0jH0r0OTvDuJ7K4qPrEeEYAgnlbV5B7Ju29LifRZ/SPnJzhzoW4HBFFV
NoJQfcK+/GTh2b2z3RJ+X/yiT+qLkIvAG/KVZsZSumkRA6hD2Wh8vLJGUaLPDzj93j0aYubh8TYD
T47J36YNdtC6OiV2QytBzFxq4eVPErfyoJAQ2+5cFYbbD60ed6xPrBbTukfXfpZANFCMdylw8RX2
CJpKOZr4YUswxlnesk72JkGGebSNSoLm7qv2zj2EBD8/lvMMthawP7nf4KjMKlz12td9joiLpMAU
FecLfTvJcFr3F9Fgmqf50tfR/ezs4X2aITxIheR0ohuOUOhdASyNzSnwMn2cGf4SmnxqC9j05wSA
nATnulN0YPbmkOoa824+TEyps1f0ejCE0maMcSR3wh8g1HECdN50BKSxkKuneUSTFBp5BeZ7OVE0
qjIMPlJwDqiwN3hdxvpmKvx9Su6IlIeDYUeOHH9fC7hRE8wWzj5dllPrDub8317Aj8KRqVti6S21
w2+578CGIbViNyvzqtSFgpeCKdEJBS4EC6WshhZnSISKBFFG3+Z9bKw+Ft/J15CcT9AHFkFAlIEN
91UpDDlgDybaeH7wuVZawl6Wvoi6iVmB69d53JxjL4zNVsdmdRfMWaopftexeagTKWbY07cqGdDY
YfUBrI7OwOJdJK2c3R979KEyqHLmWOQKJvt/WAgKNY8zMvow8hpVbjKqApBPUJk4KmrvdW5GV4tn
1+9V7DzfGOZLImIByXTJf56txb5jsMPWZE7/xR/eE5zFVeCtUXKUcWkY/00Poxxh1dOYoV6YRDbO
4lrfEUQVxik62NLT2Gvk8fHEZtpDnkUDKbaRPPJQCTvZGyrF2udo53kSSKIjdK6my+9Os74IXsqG
lNXBiwbJ0SRMGC9ge4zPBvF3JK3jzorckIyGLdTD7EN6aLYVrrvDQQvEnLH09drYtZhfxAI7gfht
Evw5Uxgo7HsjkYUu6gSZa85gXlz1USaN/Tdr0zoZzJla4XQv6fxZvhIAmZdo1/6qQjQbQKkOnE0H
HQNVcE9wfGcEuKnQFIkrUAfW6PfJI9w6iTkZ17nF3jecgRgVnzlUUMFiJ2Y5N7P+dJ02Hdg0Cwrt
uQgRswXsg3+0kA+FsVZI/0lwZwyGdXPHshfdIg09VWJTmtmpvUDv79Nyy+RwekXoglb/66MUvVh/
3RE4jlslYBk6nDHgASV+XadxyBMdWd9R0HhFgeeX5uWr1NYsCmHEsLu8bwRWhfhKmYH6FfCiafJ3
t2CFDiTtTJiGURUhqHytpJcQkIX6mKTJHq8qWFw7P0iw8OvLg6MsY2gt9Hth8+GNuuAMhwtHwpdG
7wM4+y9imZsIvmDJCXB9z5DmmnQFo/xa8ED3bjVoER15sspWDJzNjSK++t0Zg48axkqApRT3GFK2
vHVeWlE0lXy7Iq2anccv2sLpTgwr5m3XyafR1eQBOx0Kdhqz7SMpn8cHmVVUvRcjnLNJFnz92GtX
GEp5N2MU3jkRRNK93zFuAVVMyW8bJUpiRC9xIBoLUYEQr75OfJr/JWYGahcWci1Ewazg4GFPxXyh
CFuLe/C/FhCy+UtYVm0CmQbGxdQraTuGU5ueT6nWf8/eOYbZ8FijlCU21edL/hh+w4E5fR+HTT3I
0JjchAcr8ftjaRIKx45MW92TGv4STLJJI2ApjGQpSOnVhgswFA9uSFPFALD61CIVtvJo7nfWcbZv
T5sws35NPQ7rgxCZaXvxC10KlHpCpx34hvqwBfUhRmY1pNwHFwxwdxV0ZzWRNhvLGfYAvNoN9p+Q
gYv94ESjrSB89Zk5DmjAWOSKsfvBbnC+6Q6PN3I3/Gr9q23fDjXBTw+z9OGKuqNcTSdDzrEIbA5k
JjY07Dn4sHpU437vyOXwuoHImABwBrI98HoYHFrapzogcD9/HmAAnGK4RYKgjmPvj0O70pONl9qj
0aeGf7GTEt5HNqPFHZzW9XD0hg14FOIaJszK0In/7LG5QAYxfT+sPC4z2sHu7hQvSLEPHvNp1RAR
Fnh2GUlshzZUN21A5RKSTdUpQodMmRAJiLBWRE7Eps3tAq3sJ6TyZRGB8IswI/ARxhEoDmR5T8GY
mzu3/Rb2e50Zy3YOXoA+bQ3kfa93gCR4+0nQQLDadxFMOxxiIyPojwX8bFLkIo02sjfXmaVHA00I
I43CTZ1CfeW5YJ2B80zOUgAwLXtDxj0cm34hguYSwixl8b6Z41l9qBkDoWxnB418XXd3PiB6P7bQ
cvuxhMlbFmKP+HDDNP5UxpvWOUjQTlX1t6ImTXr2SluN4HpSrq4Shq/04p4IRzzEpm09q3Ebj7LS
EfqlsJ9kn7ykJ3ppvHiGq8MmUmIvSVn7Y46rMc5jRliWD3D0YrZsYwICxo9TIsHVb1Q88Zd0mkrI
T286nCG/NzYiOh6bS4hXne5LD2eyO8Ua3M7SAOkw5i0UxYYOlVXCVKFobTKpARRTFzDewIMUwIBw
J9oQu6dsQNQlARymmTkFFWesnxF1CzbvcHYfL4VXs0q4ZbgJPezRmAOoj/DKCJAn8e7/MIItVdma
ZSpWjcjIR7zAc9tdRtGRnzVMTSvztNpzx0XlegKEZUnT7dAtQJkmcXM8BmMfMjJxKgoxtcPqPR5u
Zw74g0PlwFVPYusWLYVzZSLPdALp6n4weDDkXnXh7mqvibeGCBvxgYT6hYWw5UTXxO62VMklbXSd
yvPqJ2jws3aekYF7FC0UtIJr4DCpw7Zo3WQ7eooH3NID6df9P/BaO93UbaGkOvQ8bL1gqhh/zpUx
g6qJa3I0uT1wqP21hv2oGPTMw8HRjE2+2H3Vq1YVgtHYktyAZD6B0ZQBkXHnxz58LPOXLbddvyLM
NLEM9iz/UQCPTERafUGMCIFhUIugReT+8Eg8N3jnjsnoGb5E0g54Zq0OXaXArqreQrcZiQGQPcVl
RxeUdhBJ9ZIGTvfQGf0hDaqXceEasETHCBOPmlmVoWE+tWuOGaEQvpiTRSabZ98jNnuw2et+11NW
G+ePfym4Zb+RjPJYHGM2PnpHu7b6LDukBTq4dldXONNjxWQweaPK5JECFLE03YxTDBJ036MUuoSQ
uxOT9DDwFY4X9Z3VvePJmOeWzz4+o2b/VUWTi2gncWwOSeH3y1DUGfc5nKpvAkU/rnwYX1sSdid9
5dV0kg5Ji6s+VNRXdP+Q4rGk8Sk23pjtnMTh+OdiayBfAoBPrgM5VGXi0PHHGeH2ZTqBhxvW3hVR
RcX2DCsGaueU0EoBOgRk87/7mx6oZpCxcKrwA7tyc8Bzzk2HnnGW0JQPPu+Dzl8b7X+uyuUidVwh
DAdm9MyG/WT6WWEEi9VEhZ7h1MWDtKLyvhLmFsokUlX+xAfEiydRop3rOoqnRtvOfr82KF+eRiCF
WCf0gYLLLhC6Z9LBnI96oYXB4pizn6eo8lQfiy+cBrI/PpGquK9KhkG14P6+bPVAEMVqd7q9xO5f
vgmI9fnTuKGe67P/PWpXiV1zvyKjU3GjACfgdLFvBnx+LcLBRANsVSsZvoVi0/tTuD37sSLf/hjZ
wWweSaLxWQOVq8V3JEfaZa22Ed+mSdq+ShREAy+sOa1z3ODDfXc+fq7y6A8/2/yZYXceo12prGkN
jC6W+5FNq6rU5qhE295NwPpIiUhqj1xcSnTvmol8P15AVWg7BF7Llx6Uq/T/A6A1R4AgmiFbYXg/
lUERVapU7zMJ5Y12dF+FEABU9M78dm5MAKdDjWVSMqmfLklR6/Bmb0gOmzfpcDg2rEHAJ9pSfs2K
UGVYgAGHuSWCWaLShpOr5l+wqSOSUxnq4V0c3VRFgfqPmiGs/Q7uTtwcaL2pJjvFBwumu8rzYYF5
57cQ3grnglnVCkinkfzo8P3L1JkpJPpn094pgXZ18m+R38BE8LpmNzf6OVuIA5NXXAu/r9W2DFQi
S6Z1J0ZYyxEKoa8ybouiAiL5jBeG8rTSkptkOwSbR04cVGl0XCoCzPI37Dvo2T7gAE9U3YGX6+Cl
7sW27DKPG+auXSbpFD0zPaEfoiySCrf3s9PpXFFEijId2eo7+uW2ev8t60pwQ919Nqw9kZxreCRT
5KixcQs+PXzNdlXiW5jxJ7BnSj+2yEHqIpL4qqk+tTPo5byGf2IR132m88KxyPFSRHCSTpUrqOqJ
1qSW7oc44BRYxzaDPmMmV0d9823iV6/5pRcq9UbppVPwXrZXBBwjRnSiq3e1YzBw0HqKRxawyjmL
RuPwv3uujHTDvRojb+u/0dqDLM9LTL9qLtWz097g6er5GWWkFUGw27pj3bDn2POxWwj8MxjB3flf
Lfn6gfkBqEqvMqWQyvksqB94ozNmQ/hlxOibbxFO3R8qvrH/mvadifbMS7B1xxWnEMecIpCC5CB2
jBYpgZhiPvr+TO3Ug0dChaD2ANVtfdQwt/h9QyhEEL8UrTFHOV/+HmFKcliY1a9NpKNu+fe+LIOk
rj8Eyp/r5c0grG5bLcDcZWd4f0bj5uwTSkyByOvk/f8YHxwfpRgy5GC1OUEtzW3dsn1Ojs0Kz2js
dH82uePdhKOYh3Ca3+dZDlg/pD0jsd9olICYnPPGgOsmOQC8/B8eMUT0xcaWfvNosw38jxTmZIe/
8F9qFsOwpvvpQofhL+tptNVEQaI7bPiQyBG5kiVOs7V1HJqIiY0seAEQreD525Cv9aQwPuREfwIs
kA9cX8iClzrRlX87TYxbMZ7xxnm8fWIB2JaRgPFgI2ols/ed+2HPuwwROYNx0Ikp5pHaMzdljDm1
sMi1i8oLtRDyADU86LYz6Umwx0ISrpi4G2MpWgXI/Hl1mKrqB89gcNrHEbeJIIvd/p+YabJKqk5q
mTYcQ1wVKuk6jyV0kVNJj6OfN+3PWe0ot1WsbXmRiDYjSiAkkN3kvYa/4JL3G/VkCMdBO4oxCUAw
QEqMC4iBg4DwyiuljJDnzCKNuNfmmYnK7PlRrkNTCWj/nd0QLc0RdUvlaKHU91C61RJ94uoFGIhR
r0vS2m1OItcB2HRjIjrCVmdzfuu+eZ6kiC1oZPzaJWQlX1HH0vUuQnwdg67fSu9xr/Vh68qBvw+h
W+qRef/iVWEXs48LbL/Q9KoA1XWwPAtMZ3w9BAIWRHmB0y06CY0h3e3BC/jLRioHXO9FVWhYYPQu
i1NHOmDswnfXQNvGE7ExvhX0bf2vNaqzQOwFmKE4+0IJhJKA+xJRu3A8RjJEjLQ512yd6MG+WNds
DucF5yFCi0pQoDnzMrJDI/61PCvuNURositQbiYNJWcFDhw1X6CqWsoBBZaZNdG7jIbWVG0tyzFr
V0Yez42FTK1Zfxb6Biq3H48ynIij/vYm1Ykkr4Gz4CpNgUGNqJRFCBsTBv1D60emN6z9eRmDIbyl
0esct9O4ysxLVgNOyGpVtghdpeCykjmERtLvEe6KS1UjFVLrxhFrYEjN7OVHPGV41CNOZEmTKooD
gzf7q6qBpdJZXHmczhuVMHshYY8FEBUbjNtSZ4K8p9hlEwjjTJTMBH1TGxvXJiXDpcEmpA1w4GlW
07SW70D1udU1IDAA3XDnmUI6IQRNwxT3hPsWhR6WBOHTQpQQgws73tA/pH+a77Sp9viEhbVXcHzQ
6tjbJ9ItQs50RW9T2nChfayp1h3j2t/IogRS7Yb6d8aIJ8zEaADOFr2QkRpO9V+SC/B/JKAEmKMz
qIftUhWtblNKu5yNk4tlEVlbOaTiyzWnyK3gESmkMikbSMDJsZhKD02ioRpJXqea7fsbtGrHBwae
J0DYnOLQKql/vBCBBfKvO745BQHkDZWVIIunvouiAdNTd4U/K33MgVdT7ZHno/3WYjBilV6E3LwV
SzBaVwx48tj2bhquHYng2pYOBUWKXtCqgYIHdFjsUQAXuAGDoHugewG0c5jiKDVJmJV5t+kzbWFP
Chu5ix5ddhyiu012rN0PMlHjvuz66wZZAWs+2qaglgkxtdyDPYtIPXoKkGlFVnM6SOI5X+K+lkeW
shN5f68pgI9U+X3OQe0fHpKfk35VZDTAx0D3cX0YwB3M+zd5dQlx4/qH5GiRCygc7S9dqkKJ9wJv
M7fJ2peQECoFAmEKEE232rw5pp3t1Gq6UgVc+bTaA3oMtqmDnvfIfwQm1Ev+7tIJAjJ5nOassbpI
ypraaeRtLcmkn3anSA/UrS/i2BUz8nwPZHRBcGAMHOzpDdgpAWJE3vIdOgbch2CSk/pvoaUKao+I
1Nbd0X4MmnoyiUqPgoAhx7oCL1b5JqZt5uTDtjEZ4hKsVJk7Kx2LQRl9/FJPx/3xtmFaawHJFESd
ifhkwSj7Q+EzdXlOxH2aGiwspWo373OwYhB6DiKfhSxgDb0nL3gpwyDWtxLyfl7bTwoO7voYv4uj
FWKOiNX49UhagjpQHdpKDbnLPHLf85fxMlgOuyN4FkQaFOa/3vHsjLf2xN8/HJM2NIxdiLqsn5kn
IPjf1hoX98FTZscVWQK/Kbb3FSwiViNfXXCWxtupvdpVD8OS9OZ/6L/l2oPZkC0K6Z2xpRljoL+w
//G1ZpvI/np8X9NCL2kdTFjqhMixZmj7xPnGsh9qbbkZmIta1xFNRJ2thSh2ODdjUCcc5zyyj8aa
inUXl1avlMNhRRV+9zq9nnpaHj1FibTFrv06Tt5z2UxrUtG3Oh/ooEY3oeFpXotaE1ye4beUYGb+
O0uZdXY5RYjHfBXenZGZn/YKuq18FKMqOVqpVGV9Dq+TH6ZdGa9k+zD1nP2cjPrkX9yIGtApygcs
zgokEFN46F8Y5xEnP8AWIdt7LaI3L+PYZ0a+IJ9CcgjtkFi6rdxeGEMz5Pv6MOOLBzBL+M1UaZqP
gEADC92dOOnUZl2PBmW57K2L5wmDqvHHHGM8KSuMozKSC2nhm2OilrfgktduC4BI60YiBpD9yjpZ
5VuULoYIzok1seYmjfFuaoFSEgZB2SAnRr2I+CfqWcXRk6zzI0KlROQnxhbIHYIdv3Tj72WQK/Qf
7uffcRiyIC+zCuRHy692IhB94HwUuAGaiwOU/RJl2SYVB1rPeZcZi8muT7e7hBTY56o4YK+rivu4
PxE1dAyGDJfb7aOgW2nRsoJyzGA1uJmbCpo3d08SoNcTgSqMZ5v+pfOHpBvSZOFjnffU373C2OVH
IA0lOrI8ezIEkrRu++HGySsanpoSbbjJ2jQcwVImY6IkuUYAgwveXgWorKZSjcHltC8IMnBvISgw
+lSf6R9kOz8goNvFkFVCPQ2HVPdftlYHK5h16pXpG9jcaULqAGeOQdVOk3hAHmfVHbgX5PzBe4GZ
XKbtM92j4gpYwEKxUbD0X4A8wLNqNLPPJROg+Qs83uqtzLgRaqdNQ0jV5XkkU3Yp0IAAEM0Nf4T0
kCUcK+CZ/7Dqgb2beqh2Z+7rj+n1LsDXCLJUdgGCENYOs7RVkIN0cFD+5ceFLx+zM/yxZRBFj5cn
/3KtKDMoNpxbbEZXfzVMgmXSIQUy3bFi2u1kV9pT7xZQDd0GoVhsGCWPRd716gYsE8wfWtBd2cUF
HRyfcY26KSVM3RqsEEV/IU1i5pWualP9GhjmjQqKrk4sgDrhHZA8uPWcOlQyd1r6XtcSUu5f6T/7
QHDxVZdcl8H+azNvK8WzhE5h4t0Dk3+0Oa7nu36FBkCeUDg1jYKqC9Aldt4jeRu7AlnhiXhdY31Z
CT2z599ejtKrNt+Dvfdq+zMqAnvgmaPrvXX8u82uib2oBY6stiMTWfj7GtnKV5VoWmeMQIh432Ia
6iMT7K+MFsCyJivnDWqKUkOYsRq1jM2YNOvBp82efRBLujY+0rDhZZQ0ncZy5y+ghu1w3AH3odVW
fyzegrZqmHQmdN2eGoFsJ0aBEmqHz+9eabxJSb8bB9UcB/RbPKGPFpKyePTifqsUMSe+fuSNEMZc
h7a+16xBcZkS+clyYyBuDduhi6JwM6ERti5q0xLNQ5/V+ITF4XFr5d7pT2iixjQ/xBMDwtjHLDVk
KJX4uVZlsAwAJw0x2ztG6VWfza5KE3K7zVZHjOoRRtsXJ49wlQxOE/z9r8MKQmjHWXmxhXZ0P2OU
DJi1B6GbaFjb+MhP1Jq5Z5VcsjeeM2bvkOc/of2TS4Fgs1W7BQ2gw0QsDZRRD9soaI5GPu4xu3az
WFN2gYYwExz3iXGA0e8o/BRBF2nPZf3Z4FWzTqqVzKUs6MExiwFsrdboqL1rs4CtQplJhiGueBJy
FJ+Uf5gaaDgzXB4Crq5oZihaHyv/jiZxFkxlvnMKgbfre7QTZQe5d0zhEwce3UXlR7VT3vIe0mt1
+MeLSLBKPCy5wZjy7Fk1OwipOKblSMcmdNZN3J2MTQa6JDeXnLhY5WF1wcaQwc8BuBj1EV9OORlB
qr9kPi61fi1/4mPTE59PySSzeF8pMxu5uKzm+qT4q6N4Q1GUTYbsaTF7ZhSOPv8BvDpCi6CHfqj7
J69uiuCkST9PaAuprPTsMGReOYLPpPuB25gOhcTy8MqO62GV7IwyMzL04iY2NgnwrbGwQ+k7pJj7
LvLw3iy0UOHzYSjTJ45G5+4w6Pgi00JqG4dIAzr8GPKZIywsHBLoRS2o+OzZXLlfQoLf/Cc0HoCj
M3OznhToozVvOD7Zg6a7CTYLamOJBPvf0Ut4PbCGI0yowF7MDRTwN+jao+nqaHh9uDMpUk/El6wR
sMDcdPBW/Z1RYS1XDt+foABX0G/Pv0Ru3DFLIqr2sGjgsHeoDQOY77Rxghz86d7UHTrVyPJrDPGd
13zvenIavbkDcJvqImd8jSLd/gqC3QvcXXjeHwR6qMoxhoRPvwP8p1SVfAAK29ksQs9hj25D8eRm
sWBTopAJ7505lFTO+ABcEHduucou5zzoRrQzjP5dxCaKUd0OLtN1gkNCNyxAL9P7JFJtubP6I6w8
h2EPDbr/y9GFlA+KAc47QK/vZiiilVZPdwd9Yh60J8bxyZSlT66+vWFkOWPurIwq8eXnA0tuN8sT
wg+yJbJxkcSgSMBacAUfFZ8Ma4ZO6S+bU4G2BietDNq1wZA+WTqP7JkODmEYSqodRnMquzTWdpAx
+3R81nD1vsnKcL4dnpxdNlE2XV8M4aObc92xYy/J7DrU3YTo2nbFaLDcGrPWK9B2m9J1+sh8nnZU
PjYKTn/qyjtkWTFa7y85Lt65A7yx+yaGJP2BrznfmEo18mecW167QUNnaX0Du4FsQujo6wfj/Vaa
2dEvWbLQLvNwxtpSw2Ff6eYHYLDsZl4X7vVSealTW0827DBHQ/QJ9c/Q6eAszli7niQpBIKb5Nai
SjVqk1EoSSSCxyX7+utwAqaokOVH5nYxtGK+djh3E2NUxUBoSnH1JE8nAld5F+hEpTpzKzBZGvX7
mCcDU7IsBbhqFydx/V71t21HQXWo0kInRdH7fRRHtN16/GnJMT/BxTNX/V79BsRYF3VsSoW58PjI
Jcj+I71ivR3F6pInbqqrMg7AMIAhAvIF5AUWR3WFYoqaT7u2/uSwD5i7KftRZ0Eu6dy/uQiYKbwe
Ozbur+XOcNGa05563eg3WAlYhHIvecQzkT2ZRCmS9yQpg5kTCIeLIBQC5FgKMRwBU4VWrjE73CTZ
8WY1BGm1aDo7RYSKlRSCkJuE/xtPUDywJbspNHltNKWQ1HeQlAqE0eU2hMLA2lNNp49A9Ki5mJGB
itSWXpoYcti/g3qiNdYRzuKmP3Nh5dh0mNFkcU3Zorh3W9QQ0+uLweqBfU0CMkGOjbFVizqIqR14
gvYTOUjpMrIAJerR1+evSDgJJRN8jG4hz/RclQVfM6uIRPkVmAswNS+sPp5/3zJ0EpjhSGVaeWGO
UafnyAyzajWC3kB7TnanLZJ08Fdo86qQlTpqTRAFTyQywdpbGGIcKugfkDIUqN9f/Y+uKsZ21an1
Kz76Ww0ejCdJ8mMYoz8jX9+40KHr0tcTRpvYdZ543CWkis6XuJvaPu0BEFGHsIeq15HlIU0K/svG
yXn+IAq/hsfYna6Q0rul+yX6FQK4CLkQ5Ahu70yGVs0EMLx3UHqYZMAxrgsJtoiyj1u5XNsRYsfO
TEqvdeAmAIgz8me70FDVzaetmoeUoXu9oTnEErfNmuuEK1/N175y8cHQs0rtiinx1ijYgcQh/cwz
Q24MAH7MFdOTgpNYGgMxwzxQpYxeKAK6qLpNOYNzXJ/uu5MQ7ghu8sw06H/PAC+ZE3fzkYeCO4ab
mVHz/KCBYfQlq+WOIgvO2pf4kW85xW1MF8TiPZaA6jk/YNZu6ieoGNaXuLN9DEgjtT0uM+KcfQru
Vq5G2Zv1JJPMBxnmTDNWa+zIVIAcUjwnNnbRZcwSZrsRo6wGcq2IYr5Rsj0p9KSrXkYd9sNfbXst
F1Z3p7D+Vwppq4Aw9rnL821ZH3WW7ZRqvXVd8inQV1Ca4PmQC0QTcIKZhepjzEB2QaS66Av3VYCs
JrCjwYEMQqgUJNmaJpFSprqyZjgZ1pu//Nd89L993OYBOcKPUYmaJKSQOSZ/cbgpzhoB+AmOdrcK
s40BNCHxw3IN64SOC7XwzEDyVnLzG7eeY7baplhof1iQwvJ5DXcgvcNds9OB5IyQR379210k5eWG
CClpxi9ZUP817ORBpb9Xnc5GXId6RqisOHc7d7wC553zxa8UlojUjFbYqjKVbtBknyievOPFRp0M
ZIRmEHNHhE59GBiuDYjR14VadlXpY1SaiX9bnxalLs9z0qxhuAHQ5mzv48WU4rBc2vAuB8i8b8Sy
GOxHfxNe1avhFVvDms0/eZO7vhI+dNj+/RGbJwSBNrYWEMKSat+gNpzziASDEhZabAPAjLiiNUu4
CQ/Lj0Vy4xFaORbjVxiCL9YJhfLvPk7L1Vqohp8D27BshMAVO2ojN9CMgnNEc0eBLH/UZn5w5fX4
FzNMqEX0SR7tpriInrRzwi5xbZ8QI5KotwRizKDuh0YcSg82WZXzEqc5CxO3p04IVNPmTWsmx5EK
nc1Y68d65iW7ZmB+K670Ep/EUSj6H6CPSQvIkLmHpw3yti0kGWC4I7nlPDn3OHDUwcf3WleCC+lC
8XDrRtD8NePpxak2w26rHjj4jH90vbrmi9gZ/t4OlQ6w5u+qdbaAMBS3lfW/uVpjuabsjIVyyVQa
D8ptGLB1PYgqOgsUQWQf5dkmFC2r2k8c762u7ZQBMT3QpWg4bH3qutrPZi8ZxOdQjtcGvCvD0RSY
nhiIiEtql6Umf+McYjpmizJLepvlr7T/07Tzy2VD0X5pxfQ7DJU4rVcvMBhbQyiVFbGwefUhfL5i
y0oOVAjEEHwAIgfI6HpSqpTBnhQawU5DcTj4I4fRJrmVZoBJaqouJpZrCJx/Pi3v6A28WFc6RTnU
iTVIoHjZRh8CGR5nFPf87yo+2gvVkkHOcorhvDSdezZUJA2LlN3etCE/D7kjtiR5hiwG5DhbGvn3
+aCf6j9mI/wDtiMtHBkpxGGx//e+OTDEoJT96JBgLgQkvnBe+A3vlprAXMThJfxf2acQ2ttGjkMu
1eVnu1IK0kpbYQQrru1gNQqzkXKPBn/O6WYQoRJl/SwrLmFXfh8+pm1gu8qun4ZZruXVgs2hOtjk
heyluK6nr54xLAMU6+kx7oI28zWyk2KOqzgiQBA0VDOa7LaOZyOam5Gsio14Df96qLDTULtPPjQC
mylPuJQAHVnQXC3iPdpFk4Yunm36rcCFs1/Ng+9bvIXzXcYFDwc4P8ejvT9WN8jA4AIIIsxn+Rpi
FVvO7+6CJtQVC5LSR7LD6wPhKITY/QKWF4LoyHErZiqV0SQjkGtt9DIG9NQVzAhfbZrx8+d9YvJq
pB+RMeyDJwZy3e5s3UBIkbxUSXmDXqflfqSyrFgAulD9IXu6d9jHtYsSNOYn4muzTJdhzVukglU/
Tvq3t1IS5XgeJg1ZylgK8tUIKyMN9PIsxZ52Ju+9vn6MFOnPwM5E5tkx0DV4ijqtym9+Crdr4kC+
+cm82LCWHLIlzQj+TowvEOptT2CTqiP8vJ17HJZbzEmte6v+y7riaPrZOLpyD+udsCSyNG/7SQoy
hGp8+oDtZecTCtz3SdbJSqqS2JkvWppcZLrB07H30XfMGotfZbCda05cRac6PcsnqaOmADVi/GKF
XxUfbwFYNEccp06W77yvmVihwWOnGzu5zuM9sH0jHE7j0Ql+tfme2xqgA/URha4BldXgmRfqZwg+
BpkDzIvhtolt9XbDyke0+lw1ztcfZIFb/e0ybwaq+GrgXBTXjx61YSVRBK+lL3QRQADjW5qLdgn4
iBqNflrmVvAvqRUlCdCAgQgZQYCuxmP8I1/0J/PYYUH8J0OsmKZq/N9WOlI1bM2rCpdXQVSgRpcn
v6fcQWLJmdLIFgpjEz5k7fh0ysyR3pyUSFwkKHUkFFGyKV2HnybYIsjGkxM3l5jn4G0FUofsWcJD
K8GJessIRGjccL68lGzsGapORYYo84JLNf+zUbQSC87TYS+j1Oxs4A4lNvtWSNdndvZgh+YqoJ7j
+VyeEmz9v5+GW6P44VkIhMEhMY8QCmkxczsXbMbbkKtNAx5e5ah+rJwKF+GRvuJChAFtGmM3nQPu
wHXniL1B2TpeTarj23AYZsxbIxz9kMLTWBZ0sQ/MD34v1+j5n6MzJejqCkn+boiApixXj0lKhh5P
mfAPZca39FOkaHY14T6QtgD1I2cK6s+ZVb49RJoy0OTiwjvvUWx24lIuYP9/B+jN5V3tIQwin/8t
3IqDWxPGtx7Q+aMaTJ1dwxmEh/qmb2Iv0SyohrEGDKKZk9vGQnTJvyMsuNY0K/snEiozvSzIFzz7
d0offXWZkgaUpfjMviNglm80q4pwr7kSCKptGMU/A7ApaBWjbqRCvu6OovEI4osrb/Ealt0iXeE/
0vY/E/jKHql6rA2xGZEEB30tg15CebAgdh4qb73wV/hmCme1RGixL2fKwS1fdEXijGtXqaEOW9lG
d+ytp58+cP1YXIS5uD9ew3cnCoqkqjeIFaQ3uNtgsfO/1/BL+QzTO6hbpkU+vUXY19xAgKZ8E9Y1
9z5xoe+YaPM6d6ko0/YhZylUyMZtXTD9Gvcv6TYZ/PwLQjFUPFlwO2TqlV/TjmmeaeA91on94nIa
z3jwnx5Nm3CBVE+NL0fD5mXB1PxZjt+2J2AA9aWtqfeQF1yDfZQk3k1KJgzy7p6lsRIUzLJBrzQo
tdLQG1cAXYCQ/EDaaT9znbwbUath2rhlnntmw0UyhNm0FJut844VifmrHJb2uZZ4esmAML9TlYYa
cBKIp326x66cLBGWoHbLvifpwbZPWR8FHISO/foGl6wXwRPO2hdTgtsNYYSMV10zmngIln0saCbK
pLuglje68KveHT78ktjOE3xya9PCqdS4TZCjngEj0904e6xhBbtU86fxbPt1eFxOyQTZme49FTR/
JeW9Rv/rm1UB9G3sx9LxKsfbhzsv5A6hzWQkGinduuUOZr3f4/7VzzQb0dwxvtPFOf6Jkr1w9Ob/
UKcPALSQk5wYzU8OxeByvvS4sB1FDeRLg0bDNoibK8fNqcE+HG5qCJnYfbT9CdcwSp382IlKxm8t
OlX8hZO8R4KFqTlRsr+MKLLZ9UBP/U31Hf+1kAqYTN0a7CvAuAwIcwI8tHpWmF/uSy+2UgmK21YB
KyUj0j94Qeax1ET8oE0hwYrP3GH1WjPE6uuT1XpJBsxutV4PT5CEKbCnDk9Xr/ASTSoBnSsARRzp
hlO/eFxXpj+u7YsnFkM3L+THU/A7P37d7AkaBuYCTVeY8KyXIfvVy2o4sfZPOmy8wcZOz1uMQfi3
FzmAt3Nz7FVuG4rnrV95YCiy9BpGpLFPZ9qzR/2qA/c+XxcVoSxBi0B5Y5enbEhW7Cxv2a9q2qFZ
2dQdgFNvA6wUrVMe5v0gQ5Dk56HdPcuzuTDbHvVFgv/dJICmL3h5iIkkwhH1FTRJKIJHls7ycZ1e
9Fze2Uih3EJi+TUbaCVt5ZiM6QHqjYUshVECBh2R7jflne5V//sTKBi20EHy6RISajR+WU2DMT9c
NIQwgjH8hBlbfXgU5GqfZC5m8F0Gs3lV61mHDRHlAwWF8RJPqcOketBQRE35hPEbPiqqClzTJdrr
h+tfyfEYtAxJdrualIO131sTGYlmyLb8yr0YhzKSSyIm1Sl2em6Tbjau4xJ3aaz5gbl3lsq78Zw+
KauE3drS4/8LxMN1DsEbKV+y/yRXlu2UtIfxXqAsqVVthmyI3GFHGD/7of/nJxBUmd81/xgQbtI0
Nah5Bfl2tIOTEK4jntFqbhDqZeU6H1exarns1PQhSwMUXnh10nM0lgWP6LD1dfSK4Lf5tLTqRnES
yfkXjWvUUbNS+mpVOJk+wDi8PxUV9mnyZkrAlwLp6qPfehGHx4jlE4Sk7AkQPLPPx5/VQxFt4l3P
dLp6ebRTMsfxh37O5TZnFgnV26/G2sXszW1OL7G11EArFUWjJEZYlKcg1oex2MP2UwO4/39N2edy
P3y046ECakydOs0hQDMSDoX0Kzz8bAL0X/WpWnuoYs8F5F6pwGSAL97YcqjtgbefsYzOnzUNt/uO
PWK8sEtFG74HTCVVe9gq7Q6K9bZHwywkAxIqITibr3bgIQW4oly93ebIdaNAX+J+fkuOdR0Plljs
Taye+MzAUsIAM4ffFQZWxeb7XFk05qQpHv8rolLOIxv/VK7yOBy5rl+7ji27QTR2bPmpxf2k5DHL
E/54P3if9rEneBmFjx8/YFaxQzRMTZbm5NkcTYsYgsdPtKcgFYJHMzi6Rm0vdYkfWqrR/uUWGCCy
l0spxNG0MibuXncr+KZx6j2nv1uUG3wVZHwyVJTnp6KuciFPhHw85XzPZHIKY92NrKJJWNWLa9AJ
cnkaK2SPsXKqJUhgRT8B1BYG25Tc8OhyehLaoNfySV+t7ekm47stkw/MJv9AW/4QfcN6OyAfggc8
LaBTDl/nIweiXT/R1KiVoDjLRgt7afjNvOkMI6/VJiCFTiNm6PyjgUPXyuAcRABSuj6E/47TMya4
kdFCJQW3JzK5Hg6CteEQqnqlgKiMo/K8Yh84MdEOCR8UPAFBIBJAAyFJspfHabhmJKY+jlZ9BfUV
8kSLxOfop+6jjrMJb+T/k0YV57hi1g9/8FXZqgJ6+IFjd/Jmw0Wl1xBTRlTMaT6h+ClLw7zrvEWv
1SbGTvQoaiXJWwNrTHvAHD7n6xdNiatKNiqppJSGzjG7PozvgEiXrMJpfhJUMv+YDwYhjcfyOI+c
bIv5sSS0eqbumC7WqGRvfy+9HLjtD+Nl8c40ti/vkSdcP4xfGNIuSZP4N4jNMeKbQv4xz/3YTDBc
SkFB1+p8gvHokcorMw2rJYAtEIBPUkySe+VSfmd72/FPCtRcq880VRoboyBec5CSGItNrleuezlU
v1AvVAtsVqq7LM1coKYLmfbWDDti13s8QAIPFqkUbmI3I5MDelLmX5zJBoOuY+0+3dVQZTcn6V8N
4mWlJPCQB5npnoRd17skI55Gw1jMDRjcD5Fj9soVQ0tYO8sSaY/Kd/tJkJdRDgsAri8F0d5I8625
ISnaHVPas98hrkuNn2oGgiS+wZ2n+BuEjJcKCs7sOL3H82kT2Phu5I8wh146c91pQ/qahhmHjkt3
f91XREsZ2nlGKDrkEUehAnO7gSvgR6/2ITOJggjAHSF08ANDGK4fbBC6aLDpszG1Kx+Lc0BctgVF
XumqyBrxp1mufhE9SxJ48bpj18Hq8t+UXnMy+ajPPUyjs/o9j1Subk+0D5JKBn+uMhoatnZwAV+L
YcKnUoZ8XWZ0ur3nAe8OxzLNKv0X2DVWDNRqi42fYbuIMrPaWWoAK+rM7FWQMM16ySRvTRFDL5Ci
7cUw+utByfLzaucMVzdVZqa0qCByY2I8rW0MMqF4gnsLrF3dzu9yVtgYE7PcEwChq8eLZIl/8ORN
a2FKrcWrjDd4O3gqR9mtiUCZC7yQSGAM02EfKUDVQzxtx7AdsGxaF9aIxuvzylFLrdrNE21n1Qxf
ocNgJOFoLRwQbg6EYgB20HYtQ7yTvYU7obYvXlAydKAUTFYKu5Xn6EDvuk8ld2yCC+9paj1WXkVO
mDNcc2pOCGYIdLax5gBYqvSif5/LQWQMz7BOlTGjQ/FHbRW2vCXns1/dX6/MISuWSh6xEbs50BFp
uMEic4BJkjGtyPI1Nly/9jzTD5PciFd+hEIQtfgqVjbAYeJCszyuzeuahvwr4XH6XyJd7whmizHv
AH/59rYb5ZtMacpCiZFzw4Zz9n/84WlSMVCqnbeCwpHZODtYC5S1Q67CGQVt76xJbSAzo0rOEPNJ
p3c2PqpKnTVa7xPySzW0hen3nth68TuQ2CwWdOVFD2sPan7NMHBuo1a7zQfQ8BjnVP0FGeZ0o+zm
Q8zuSdxQ+58qKxR0jp4BibhLonRCiJfjCZpdRdWOk7MJJj/aAEEb/VFh/StKu35LswaIyEzNs4fE
Ufbt9dg+aj2ScRzkD/SrGL0QrH5wAIK2pMDXya210DOxjktaZUj5uYlnhG1hw6v3v1tPZf3pkZDc
sxcyUH2TvRRx6TuHegSDDm+PmWk5tDHWs7eUppH9FesftJ/Eog1IHbhNUbzFUWdiO1ilyWasMEpx
liMtCge9IamNGon+/MH2zRBbLR64xC4wQaldlgKUGJDzOuHRqQcyqJE1zbXjiXBOnEOgcgXEQ7op
QmnBtlb2uHPvfJcBYMm4gxLhW6RRt0X3WrDKPsyR0pFcAEzABO7dsgb/9aXB7HiWphGctJ3Sm0eY
msP304y3iMaAG15tMfQgZfR/NorP4fTT9hrktnb+LKtxBGHeZwwy6O7tHl8jAQremGQEi069EGOV
R5o2HjSNpFyqLfr68FSZYE3R9RcUt8fEOgE3Q0r1zrm67Dd9/Ki2ArPlvnrWGXwGbIGQEedfGzTV
uDrf4AGdw0G7LG+7D5vCDyX5+WMsptSAA7OIUirYcoBxYaSur8p+Gyg14ZxsZe8LRDbkG+tg12G8
Duv6qQJ5uy+U3DIgXyktpYC1OvPM/qOliHiOdQ8LGehmnmFtwq2ghKaqFMiEUeJKWLavE7AEBv35
Ja3FHSp/tCBdEfu1hn2bB26gZTLbp8Lnj2xdhkRLMZYl2lR6zXKIfsJHqC+kzRJZYlQPK/0e7m2z
WTQ6n6ndvb46+c7WXOBxt24YoEX9Uz9z26d9pNrFfyovJt6weVPvnVl+RzDWwHzV7WAQ8kJRA6Wq
0zxscskxSkgESCiZ92HmyrRCENbABeJL48iWPS6/2Q9IshbPPjZiPlXMZu67iAjrxHXcmjIwvbph
EdnxXxoGTdeGABduQWI5O2tjtCiCjy32mDu8BdwPyQtyRWD9PJ5NPEAbaOyNSoPfZlERf0JZylnK
+ZMVI6jMvDUXhlDTIelyXcvaXsfLktK4dOaCvuMuKXsV2xKHk6pRtGSACkLH3eWRQoU2hZcdIzgG
amntDH62p2Zzvdog9NUCMM+8kwYhojjjrB2OHW5NrFgUws6lsjwxMMg+oJTK9C2NEhyEY7z6G2ut
nIR/GM2dfVCq6BSfnDpBfDcqZ/VaH9C3wZOBIiE4GSODwUcEY8AkC+RG1bWDYQNOKqAuEVi760EL
rSIx/+8FqTM7sndnUF0lv0b03JKTsmLX0V3aT6o2RHU/9L6yAyFF5on18sFtbQiLK0WtpeQQ/isx
/Vcc58quMfaihBMQR9rp2hf500915LzY1NAdyMO9VZ4vqDidQstau896yHy0JRMWKMcPW/zFuaZf
wmkGnHUqBACIq63JsyJGQYo+K9MzqFerrwf/zwq0q+EFnQw+kFRjq/Ts5KDWCiCeTFR48uZW6Zld
U7YI7BcdMRCPE0EUVS6iSmAIL8DT92eOsK4IGbZXMEla1qgNGDSgyelqy+osqJvm6n2UYOvnq6Wd
X1USv1Ej5Gnxed/mKQIsST+08Kji9GHXgeBLcto1r7lJVSfdEWvyA/4i7b6uEmQeZARx4FdeQXCE
4DzFbWApfMj9KzkZXDj10Y+aw++iMt0eZ4qnEqez8yLJ529faGC2AJ+1k0WZbenJVMJMfDf1BebR
pcmZ92JNYUVxR6bPaKpqEz6pLv6phbUlPXjWcLarTRvCUQZSGda3yWBSQogFBhVOzEsdlt67uGgh
9/C+C/5akBbHhCesB1pj+q2Xmg7Nc5z+65uNTh9jflJQgi9IB9BoaDHbM5PnYQK9UluM2Y0Hai9r
TKokK+LiLXnsz7BXdXo/gW8wiJjUgbMsWnGmisxgImnw8aHhXs+awF6hGW9jzveGAjltXicORZ1b
clj7uSsxR/pEL5L4lKClxHoSHl1XpnEE/cHHEc91ttNoxzEYDiEnUl0k1Wwj0N1SSf0hwvmisXaP
L8bGOX+xScEEBXn8FnJJVFpjaUG/d5zV5BowSTr/mQAUIarrTkui/YXDUy9oMchSf+NiTJiX8mLF
Tk1ZI5i8K1IBeFTTayBAGd9eq2UNVcfyDKschw2ddErelKvWW3DNmv6ddP7vAu7hS2GkKW6Ugmgi
J/C9qRtV/mOPmk98zHPf64cDVUrIMt379xOgfK2En2oy3pzVdZf6pFuIWYg5EkVa5fbSTbkJN0nf
pwnk8fOd3o52+J0LXCA1SlIU8Usj8qAMAWwvToBSEAGMFWP7fdgqDyTEzR77jiWzyR570vQH/WBZ
z8dens4nBrOfbdfceWw9FL5kN9h9ysRo9s0+cq7V5uHhTd24lP0sHRp/kwR8BBd7OsQbVYPebSy0
NDkIaOM4tfQU6lP9oN5oigKU/NnT7qDS6q/AoUcLv9OdBQVdbO6Wdl9vxHTQw7+LUkAeTeN/a2dp
ZnAXOvk7PQvblNYCo761IdbAezcqz6NmUuqFVqH02AAa5DWGB9ntd6C/n9M18IQl/Sic0UTqAYwO
EUVV3w0lfZTbdvwzA/HTjXb4jVzSoB2S0lyco/Lphvg/vSUjClqHOoBLaSUq5l8bcNT1+neHfXh/
Gscejka/HWCo6cm9QN1sxCrLMNtp3jiex/Zs8xZFMPbE0c9IJh97QAFY4sWPtOdoZxjfO7bEIw1i
RZwaUALMji4wddce4D1ihA2yqN8b+sDkMHL1l34H92Ie5nMKle1Jap+nvkOYrFvtoSsiO4h3edwd
jVYugqzJULls9SNlnDv5cnqHDZpiR/KfjUuhKxu6qUakRaLwa++nm4BKxEjkdKP4kNL8vDUNJBIJ
iKFeINUekkfPo/qzPPIjSytGyuIrWpIXbIBClQmUxQSenQIlNlHrOVlAlGO1+MzXaOuJeoW9DIk1
rFLWxHdInoV/90mw9HoSBQlSaa6DzGv9Ep9GCCpnudp+53OA7yjAnQq4bGxuhedL1wRi4F35iguh
RNQsV9ifOAjkcklg23ypEN5mpwou0/9xqzNdTgpS62SaFvdpw+axgJb1z1S/d5LdGjRfJOzcXDZv
V3hBjFASMDTffpN6+kIzbNxdgvLxdDkQRDncLfjnrkUsir54iVC2xJvQhGQ5xGQp1SMAOF+5s5tb
QhY3zEcomIi7YdVx4H8dUrFklSEuLzxmP7v1ItoZ3JT+XOSIjQibGGkIeTD7aIQsVk/iAduhjOb9
wSpDafUTsHYpq9G4DasIutShtA1n98pMpZ2W/mWCycv517fjTViD3Nsl3JuuNgEWo09vo94k2Zyq
fid4bfN/I4TSJOhde7dAcezhk8G0wHJDebnGjbBPRotc0P0mJqxDoHc9DKccJLQn+dW5wPo0Dcf+
kL+U7wA5eU7CzAkWkVQrT9EF0QiItHV5+G7ozchcSxr5ukDWdq1HIlyr6lSFSEMMGiQF2R/bhWQG
o0576y5tq5iDv/GKANypFl7VzQaIRe5CWb/FSfhR9jJYlA5uhS9JBk93iJNqaCvAY9igmGDOs0S6
MAfi5oYMzoLwpIpRLFJSfW925O0RlQCLP3C8o8bCx24PcwYs36CmjC+eCoY53zG1yv7BrqIjRBHp
dFtitryO2n38l42fGhpAJhrl6AxkfIZDI2miIkgYyqus+ayfeGfGt+WEAt3yCKxKCZS+hZOvjl1N
9GPhkecFTd609BYvcxXgi0AdXUQ/zHPJrt1UxCHj5LNKp86ao4Ka+JnKOS+PCGBxfIk+Xr5WnCKv
HA8mw03Etw4sar2E0x9TYAU7cykEa+U/gVlg9oKLb4wSoQRtC1An5cdk9VAFfNs+sA01KOgux7/D
beiMsCUuvCrZZ7SBhR2YGor0hW3i9EC9AKD5dq4Wix/7GUgy3m4olK7dO3TJfdG13IxQURX4dbzj
8uvw3LSRuine2cqXqPErll+GStV3vL35+WkXta2AHr77pgv6s0T9s+HtHrpEAQURUBn3jLr2TYYY
WaPs3MhJ26UamDodBeFpXvdyloVUGGkidbAtrj4LfILbL2DneggJDMo1jvOsJS4gH+dPTtx9+sDx
zdSuHSwc4l6Qfqx1Kh+mdvTQn4DLhttFeMK5osdqJisNfhspJbtll2eC0x4DmF8MNBCXJAcZZg/p
v7nSa1c7wpJzx8jAkEcCtcvpsUbxhNoZGqYEkGFqagzi6zgVVCYQ9d6eMu6bL1LcOb54vWoz7DNH
b0Z3c0y3GhA3+/sdb+34pG03+ACp/kUDDXFp7mU8b8FN6/OZhCuc3WtVsxC06Wb5sqnBPP/DUKQK
U2w5dr2R7mGVjnAWIHamYxHqP9YggIZPf6fJxAleQo1U/ueybN2icK7Q0qF5fC3j0hSoVY28/7DJ
V1tcHDrQ2sr1/Qe6cwqafGRYex1hmXOv8dCA+Kudwa4wVPOKzqHDYT7TybzI45y2PsYgVc7UOcvo
zb7ezCTeg/tUMnHT+DTwtonDWnZ6oBUnDlCNX2ZNbPBus4Zsv780ufL1V+FN4O8xpCTZ1cEjwS0p
MDIiQyIt22Os7fbVcKMHsMC+ImJQqCWU6Dm6Txb6uN0joFCS+MpntFb+Y4Hd0BtmeFtnSUUSPoKa
TCbt2WAGQebgdaODYK9Qq/AdqCofG442cZafs/n7bv96VorrjvK+kHjGnbZ2rPqIQ4iYCQCYh9SC
fRVaJuGdkUJkWHXaM9FFLwVcrzUGiSxXXI9fVvERbKPt0yGSP39Mqq+/88xea1lEXqQcx3Hu2U3C
4k897jPaIK6yCTnD47ZWJPRgoBGZcsB+pyWzQHmBmq+ZYZy7l3aACh6ibGYWXX6qbHbIJnMqfQjr
Zp+KnBBhmzzAVNkVxI5iIFpX2OApqpvAo8JrdRVS79PUioEWoQ7W0GGpVAaJtHBPN8oGcGCeSys1
s5Fkz7JUROTEV9XbzfYeV/HK7kC1I+wgfad3akxdU0l1IaNdXcEK3Os06Gah80cURKac4XlLicJ5
ArDvI0lXvDdWwvmwX8yBvAp2H+pk46OjVZdMEd845l1EfdoIWbTdd1AUnnXc4TRbfBlatShJVVGL
3ao4lU3w/eGTUsKmETFZvRisnTcUCwed4/X/S3N3xQlCQz+8xP3vEbTwl69DXSJPG3gDQxkylyZ1
sBDx0uLV+65jbnCcEyo0RKsFEso6WC26xHUGkPbL3cwgFMIEGaHbsKFC48d+Xz9Wrq2YBsD9iKvS
hYD8ST3Ev3uCSjWgou8L5h0JffifsT3STg+ekWiTPiZbcUvGDvfSShDjnLl7eJNaGI+AMRNEz4T2
ugwizdHJ+8MoNc2GqkJHqJTykjBpCIIW5cLSNxoTflQiyJdyzbb9pzmtRGCSscRh7acAJCQhMh+Y
+jR4F1B8X1+TvxamM0N/j7L/cuzrK8jNkVIsqHI/8Om8w+4g5sBNIfB0OE84uFL4tuTqOOAjW7u8
KNdubWKat7M5LVomv7bi9+XBA2ZrAk+veRXfEiRSLlRRc6Mon64l1Izy69R190zLr83P0su77Yoy
HuMlc/P3GtGteX0O/U0QVd/LpHUEcJZXRpxEuLptebvTvrZHNgpvYR6j6OeTomyid0fC00j1Z76M
5kBmANYRg3C81cTc+OLyCi4SmR0ROQbmSv767jfkWT2PI5QyJzyBdI2MN4yMyGhgAGI6cxoUsA/m
+SZ+v4Ao6pdxClc332icWYfmoyGfVrtrRMCuvOFuOl9KA22F4ZZ/vPlnj/ng/3/6AJTJqdbugjKt
g3XijHCX04Ok5PIPyZ8IHirArTakP3ImxjTMhROnSWkuljS3YUBbbgMe6Tned5wJuT8xJoCDeaok
Cph1HnVHCJNngbxmz4QunJCu7irnat8qkomJsUWPa2bZBskHZynZQa3Bgz1NDNqsu1iNjQjRUqgs
pPCka0sAOlo5V9VvUFqa1uwJslBK7/cQK0yPlXHd6kqVnMu/eH3SAcd/S70gdoBHYzy30745RXhO
npvylXwjLd/HxRS+s9/Y9UpAezj61FonbSmmG2HQzcJSwg26fIs0rhhe11Nh1qMq/TPpvxB1Hh3Y
UYmPecloGWmWbxeXs7Bsb3br1dCIK9oIUlJLVSolprSoBjueESAoej7fzAS9IbyT7uSFnZrTlMvu
3MQfZcA8lYPPMNZLnQTQt/75XgLYwTXtLUmlgMXmm/CH8JdqwA/k4i7+1IqqkQ+ck+xrTUuwNZKV
Wz+a3HACK+gC49BBBNqUQM7L1/MyXM7Sn2f8HKURZdF0cvMdC1o/8eudwA6aVGrG0gK1p1+nYFQ6
ZrVS4FtiUB0znC64t5reZGjJjdNLs0UpbhRpr8W5oHznZNuTk3wq4Z6U9RhaPblGvC8iM6PWPFkd
94/u08wP9oXG3sY78SMUhpx8iWyvos7yNJNSRBfojjcD6w3F7/m6lj1HTrHA3Vt4MJWIK/JEc6Hp
r4E+XV1NG74FbFOL6/EMD3R8YzU+ZGipvoGGKVQT5vamXQ/IvAEuO38JKblMRInmK7MC7YeFWiyj
R3hfEOQUg/ZJ0p5wM9nMxVpPGKh6e2+o6L4Pkk7PAKlx7JxOQqmv5lTFlFPIXA1eF/+LjTNdPc7w
rMLooaz2OWjD4XHujcPXcMmbhvAeOulTsEykVVHDBxgRz+VgXlPVdbIO2HbABaI4+2k8kpaA6fU0
7882juRLpEAg1DqAUmdje/ywcQqLLEKr+1iDXg6EnronfIK3/3UXoyh9M2g4TLGnHBkYWLdkNTDW
HXLjiDE/WD7myS/Oor/uO3JCW9mA+9vMH9PH+BQraeAhLm9Y8PYKPzBP9xudRGX1jHEvFhXkmwi+
fMh/86WtvNCzqlCqymca6orhYZRut+2Qce54bXIl0cq1ITLANsaN4v5XILAfXZOm+QYS/hdxeA05
+5hnuVdwllkGMu0gGh3yY2BHu+SEabccH7T1n/E4kzsbj4g8xFS5uZ0Ps++jG8P+kxyLcedZe5Hk
yRCExHVNbAeYL2Rpndum8ounMUlQJjBxSo39ScN3n4sLCr1qOcscdwMeTaL6HxiMrVCvdVzBPytG
7DU8D4XWP614Tb5Csh90BP6SQJpeZhYo7pqHIFc/DWAWqjJFqpJhrFeorAtBjI7o+uz/5P1ZSiLP
ojlMak5RzE+59wMjVoC+bYgzaLK4FIdmSmArVDAdhuPCiLTzwAxdM+sPUCPTpfNoiZ2+Huur7oP5
l3UAMjaz8IwIN/mh/8Ls+YuKVgXi/Fx4/XahxbVokVJ47a2OupJPkPFrdmeTjTQT5G5TrVYUWgNP
nzv39Iv8N5YsvOs/FeCTqhhy/WtDVb+DkBcCOi4bkXnZkNuu6bT+JnJq9EgtRq1XolotovO8RQms
j+Gg5usk6swV5zFarV4kYyNTfwPSZ2FTf8hxdMtYjy/fBS/bcazvi3GT6bmcoPaZz8ZK0wvqCNpy
ZY8MFhGoPC5/rlrwQDj6GdDsHZdAQPjx/D+9lH8MsZwWW2fxZji+hO+NB7xjCzEpjI96mRl4gzEu
a9sITjCbi1zUrQALbRXnMIG6g9CRjCh4oJw6V01raEAPQYg1MugQPhvWVUZtOigx68Z+qwq00t/l
GMN+OeQzXZ8bM1OstVbjT4a5NdXRLGQ5kdJ82aIsGmVDAtbmk+ILp/6DWd80fFipG42dVnJ5+bJ8
S+6gCDecZSg2ZA5rJPySu5j+nk4wGjSU5zgX5W9KqdlOnwt9VhzDMH/a6zWDcoS0vODVdob2Hqgu
TBXWx+4zMwj1BGZmaVPH0XoV9Yk4kj9M0LUE49Hg6cmj9aAASmWjzmkDLAhQe9l4Q18LCqeyvBVG
wHTAW4DBXBA/zL0nuU7QqposSdi8r2luOM/p8YdqWfJssQKnQUuWh7GKAz2otqXPKFyk7zMgFwvk
A0KOyFNf1sp4COqG07pBA7xUjwpyAzRBlUuZYDdFQ2d5kSyVfxFXEZzvqK6kysxp2igC+Zl/rEVw
krOfsqzcAXKWOKMGDoL52/+seLzk7cMn/NyahhG1YHM11ic5ZNwsVQBLIY0/MjuJjRAKLwwoS6rI
lzUEICyUYNYtuJEfKLvPwL6YWfPAVh69LrYnRYZeDALSgl6hkb4dzxVW1XSMmvolG81WWmdjaUfq
FB1RSLbOrfeYMo4k5jHyEoBkq9h2Eo9SB2XehHKWgfgXKED4ihEjCWdT/b9vjj+RELt0JkXhx6wl
Sx88QFhjEQWDZK8ZjscMgQFo7fRuef/YB+XTaU3XH/fUZbL9L2Qt2MCYoKsBcXbmIz+OXRjl4ZnY
Q9pm1bNMnx9PX0WBXTYFGhAlMAurJ7cOliomqZTFbnsVCGD8SmouVtZ1dFdck7OISkM4CbW1VyHc
UsxZOhJilNPuMFCGpIcNgMPiAHh45YD/z9JCeMP8bEcxaBjiUw9FRUX60x0otqPh+Aoqlob448BD
+4yGwpxHa2cCc7iXMvFAX155YT07uovW5S7bpN4XP3Qo42GUi4scFWQV2LDjvGECp/XANy8eJvkS
KW4bpPiN9GeHEyEPgpOF9B2uiYyexU5Y+yc/WcHkOCB3UNd3qkHk0gsXvcZ3RbO1cR0auA8bLfQd
mbmLJnlLAlcXHi5PF1qp7T74BbM7SkipYsoLUNhEjqN7+kUUUsWfAvYL5eGnUdXamsN9RNe4XLMB
5zkdTk5BhHE1YM9A90zLZ0FlSzC9Wja4yrpg8TURwUBUNLC8/m6JXLNKVBqJOUD31QzE0kWt3XYv
RSyJ9JRIqGucKFrMyaPDzytceMAULjHTdtBRniuGl/FBbtzXOqYtkrlI6r8nE439Oce31E+BQIq7
gkBccl3fPHFABDkm87L0wv34yhQHF3Q4Oo0tnIe9S2h24e12pXIIEUhlrDb1P43TIgemCVbKYhbI
nezkXuDDpXP34ogJ8gcZ3pyjIT8tPwunPPz/zvygjc1sFDSDkX9PIoUJI6cx1ISG3dZX+3UnrUUy
PLDuwlfV7MJm+ephH6u4+xr3x6wdPE7ixihF5yqGLmrCSp5BYzepK0Ja26R/DLO6piP2foc91KNB
83ktQYMkxVH8iRkkN6OekTGFVzfQM4MuRYiuB7ZfqRGkZQjVlXJisRuIoB7ASnzD7mWzKhWHUyzy
/j4LdaejcK+DSZ37qeMqkb2cQulDYO4E/VQsaKCtzzdXSCmJq+6RsQC8E2CDE4TFTaCdMnZgVGRa
gJ6iMng+myF+G82XzSsSnQ/hSHXXldvbzCr9Sq3UKkorpo1YFU5z3Yco3ShWGMPqCpPv9pis3iN3
N0kLgLjHsNNbbM3MQc50UjUgSB3ZnJP4Qc/tc5rLyBVgt+yFbyfexT9TA4VyTXFv18KiSe4CGPcs
lg75Nlh9Q7vzkkFJ6kqAHBC5kvb1ER5OTHVc9PdNaEbMXe3ICb1EcIhA0/K526zbTWy1QcOD0eoS
i+q+SOtXcSwdTYpKgh6TlZWS+txn1hQVaTV1CgjaHofpEau3lz4dEjMXlLZRx8+ARSq6EezjYXYc
QH63V17WwQzPqbsowvFswENwV+VZF7DyZTzlPCstQjW7biEuMUy7qjyQUHZHYQMGC8wHr5rRDejO
xGwa3dd7s1P4rJtovGZocDQU9uPg2h2PJn+Uzs9FVZMvUcNi5Z+CGq1beBuPwY05aCQ1Grh0fHFS
Lqr/DOJ1H4UAavhw5+ZG4slSv1SCbdl64/jdio6mxY0FqTom2RS3lggklZwTSCcobhxWK6GHLhd4
EmBId/zihHDeH+CI2vdc0OJxcwXdykwEfrV81P0Dd1CILWdHgmdxRlR+N0utTehom9zd6og3V/zF
Y/znQpVM0Q5XERFxbBtLC8WbNTevld//jjSVRe2svdi62HYQGtOCyWrrv7i8iQ1FF5nUJByraCXm
GAcuKzqHXMSc8hGXjdJVADuSSwblIpSWcpOxj2G1wHWioHWO+eix7o8zl4nz1vCxkngt01qDtcfr
fgWjcn8Ku8eJC4zbkW9TAcihhQQmf8dOlVv6tymXi6KUtRhNDqolMhmwAyhWG2BHcyAEco5KTbX9
1MUwsRKkTKlJS/8Mw8XLe7dUHrUWAvtpl4ALvNILVA33V9KsKANvytTmoLAm1SF6vvdD7+LJMeLe
2c00LW+90iI0LS47PNkbLrplPzXgzLozfrZmX02WaelaY4DPQnnY3XW+jWVE86dJ7jYhriASsI51
GkXaLWGl1rUbhwNoMgbszes9bGiJCl2QDktoXxvGNnn8sDpgaA5GEUog9Ps9aTYbi4ElGJBEv4T+
5hj2r7G8eaOelbd7+x4zdroOuiK5zTP3gWSAhjDDUL3K7R9uEJEb6f9BhcbId1x/rvA677pRkzFu
8C/tmgiF66xjaWkwCSY8II+aKGFzL8wnlkP4tpJ47BhgjRN8ndeKY0nIIq3fSuzZW5UEirO7T0rY
nBdPdhOhfNE5UXqiQta9tc0/dsgL9/CbR1RGv430kbNEdl030O3riIUco912xP3wbwc07CZhn8SZ
S5pMTemupyybhjHcDWf+Ggz2oHEyOpE8GVoCeCgJ6TNp7fnxtxooF+Sxi3CmQ72PxFkHWp86tIaM
j/C/WNxXzG5NYa64wETvcFvXeSUx5Ql7Bxb3Dt9tOzZEkqrGQ9hD4qUP/MFIyg1yz5JmHvuxaW+5
YfkayvqOJwrK/QAXK1h4ssWL1S6M1+YXm03tZ12L42PLBMHblHvoJG3mMQ5fJ4axPHPQbUXyA9zQ
cC0e5DGke+mWrwWfM4A1kOzmsTTMe56Z5YMmFUPF/zG0DjGpC1C0TadQbKJP3J2hTa6DrlK48Sc7
DzVPa/K58am2bJu/y+rAqy+8tRDsAaFY/UnZ3NGl1TPOjoq7kpBepD9HM+C/PrBISLVs7JVIlU6G
Evd64fepsZzo/bHvOgTJbvGUDLR5VsbexsWEcG/FrG/m/kE6u3OjcpNtg5iXSBA7baRo2D7r5jTM
aEi+IvBBxvtSdoBKaukrmVxQK4h4uEI/7XmBe7aG+1VT/0dJIa//dM96cSF1qQzJ7nhkQZHCxmlz
k5aNhOsbuMtrtiTnJtkQiHF3KnjK8BDuBXJYOq1oD8cQfGVv7tiXS8KOsip/VuUNCsKFTGmUr7SK
NWIVD10saL3BoxF9CRnwZk07NKe+3BNWi9cRUNnuHMSkxVYTGfhOSguQGbaFoZvoJVYhyX9sBTON
uTJuYQWe9kh02t9fyhypg64o+kjRv8vR1w5WCHHj+CEnDwcXF6z9Z7Dz/s0a2uKj4Q7YxIeOdUML
x/XEEEdkSVdF5MuUvcSenTlF+treMD4gmdKWnCpB7ydKOGZ0xJF0urnv1pXIyPAhebm6mwDuFDLR
YxRKRyzon1UMrGpvKZn1T7K8fOAMbgkh8v8P6yoyc6XUnc/Xbmm4v21KHCEfQfSOW2GVXkxxu5f/
Dj4+qNdVZ+3Dut+aDyD9hXEe8oLsR/q4riP+Z4TJ/RO3zmtpfLJZi5BYKaIbGsGtTQB01/rfUTek
9UsGsfbUZbWB/YvMj9VUJc0boV/CQgub+zHQ+5RQmh2f2WAOg2pdR3MqsmNlA2aSiRpwYur+S9Pi
/jX3+FAqIDmSqt398es5NDZ+9+Jjwb6th05ywHjFmDmf1LD7qs+jofeqRPnHC191Nmvu6yOs3MMq
goQ7NJ0y7dzICVZpa/SY0/mBtBNpZnEJ/sau9oqKs/PAlEb5AUWlRckBn59e7Z3MJizMJZsq2v7K
mTzonUwxDLhPQ0UEgn6BJwG9VQABSjdRsxZXwiN/2uVAWkRWIQhzUyTQDW/GoiloapmQorYXjiQK
L4j4i0SdpgxSqrYzvbvfZwzhSPfeTu7UZZd00d2o8HS+Wn434JIcHf/4nd0K93lndp3fck+gxnNF
PQfGZW+fjrugTHb4EL9/qhFMFICOftuqr/YG/WJENPtf98Ok2xo0GK0AvxhaI2VVCWcoX/DNBQZC
JQ4+LpoMpsrUOiUJQ407GrFbmqYGiv1vJL5tGf95XoNyElV8EK4+ScmcOJZy2Up+JWniplbWKoqx
W7+9n0QyHPUIKv8tg3MVXUi8Q80RxJEoDeGuz2WS9lVt5WZSi3yIcJVkIpCjrjv2J2PdQmobmLll
vziwmnSPssKSIJ98it4pFTem1s27II9jSFI11ZopyoHCo0xvwkdp67O3fGPsVU/57QeuOZo4zqnr
maerTEK5MSXJ6lBtlsAhQ5IZRayn+wYcafpmgAMZWjYP6itfE6rp10Sa471LKzhHEJJ0eHNIdPFz
TyE95QJfvVzb6szglpXzlmMxuzZhfCdWryPLZdSbz0JaHxZYLR6xR1PJ+7DPKVb1yra3FgvmoB3v
fTtNhu5CbpqAyYJP5cc1OxrkWMXbhOiSbo40CEfgESpC69gOaZ4jiYuw8sq77EwqYFPgKwZcD0hA
FwwX9yjP+1pVYgiGLENPVIlIcMyDO0vlPGPtZNzxG9pn4Tpv1v17cmljDwmiwqAx6ze1HXoXDEPT
W2pU7aO0i0o2VLTl1qkNC2bSuVSVMYQCUg0uz2d0MLyhtaS2R135Vrg24Zbk21SvFxMnlreVX2J5
QYCqxN0OaTQ8ZhpcNN69CIVSqpUstxb+vQbvmMB/mVQgvzGWvAULQtfnvfv5YjEYkQMg/eCmXHhC
AEjgZMHzjR1mSwlC4mEiQPY5+3bymbOVQrb7+o5vdg28g9AvwRyAqB5Gr0iclh7wN8pEha8FLh/w
SUVKd2FqbNrVgASx/E19qXFmbrsL9RwwB6IO0maWm7kYGL4Iqy8vBrea/3yRfid2ptIGFsfQbimW
YNtkQxWHsJdMT8KeW2/bfhD9SRjdHD/kHFR785PCCMYgihvPIyZRJ5eoWrsrK6mObWQewDnaMPgh
dyZ/hyKucxpHJtSyej/zyc6jlLD6uQ7pL3P8hfoJQJl2BsykYPbswIOgvXrSrUbEvB4XHB5XKFdb
0ga0zpFXiZ0lE3OxNC9z0w5cBrpRbfEuWmBUG2uAo/jDtoIwmawGswjxyNWk563KOdaqLVA0qq0R
gGUYt60j4ij4CWTfxy4HBURvYiRpkWZezZbGyZAQyge2kLZ5zREucnp249usmNFaqYaKNGTHqqcq
Omz53XReydvJ42lCoQNv85oK26WeY1XGEEVl8Q68eWiBI57DpD7nStla1BvBSTe5BtuFa1P2RspT
FXEddCGUJ+PSXx3t0qFfaxM0z490cRk2Ishrg3TqiIpS16KaOp19SBn3WVfIY/g/L9Fa1Rmn8Ugp
Psy8YSrA2PmZcxUR+eRtweCARAhWMRgxdc3lAZhO8VYoKKxDSFx1tDq+MAJ6CGgAAd0qe83KJr6d
fqUV3jcdgHkyt/YRlAmsRO2Bi4nZYSqk8t6E7G8DhF4jpJ2D7MO6PYe5Io0HCEWWoNGXFpReV5rp
VVQ4fLzSdQ+r/7VPAEe+85jEXV75PkOwXV0KpejhkDc8y8v/hPd5OjHW7zBjQMIWfmLzxcr2YThe
U50RR9fNyadrfcw8dlx0EwkI+Q/Fam+7RaE0vCjjuwrtmlmjgSA8Ao41h0mCRo17xEXkD2+gzwnX
NuJc0I0Lo3gCYY+pw3ZGea5VDsONl/1JMKFiDVzBE8pB4lKEYQpx9vhesDh4I1n3bV3JeRE/dTuj
g/0AC+7csx0yrdHSvlNz+dkfIj3+WX4XNXY4u2X8Fr9ju2/uCirsCmNsGI2GOEyj5fyg38vsNxvp
0Cv07wan6LvxpxrC5mZQUJxSX0SF/PFtNmxQq/tMxiLVpkdmLI54224AARnDXu6QWKcgrfcM5qWW
YkUkyeiJYx0ZdamNhBTPckjauPEJo+p8yVuSs270UrzIM0a3iaZ9yIvhNM5fgBGmZupmCOrlMBND
XPk2cDVN+umR0UPFOwyAAeIg5Bosm0Co33G6Ny6HKQzYKP7A5eD75kpv+jMCmpW9JEmr2FKKNmxb
2jcFRlHEQTX2cRg7ySxSvFxo4nX27b8NFMI9tg60BKzrA/kf4jjagvBVuelU24uQrMel/poA3l/G
oeQpk3VIsmic+qLFWfoFj/QBfpRfRXaiWhg+2lPLWvzfbE1Edscam9/eN4esQB9hVBPG27gBG3yd
LtYvotMvwCsezdV+mLLhDjIqLJP7AL4BqDBgchDfPuPGqxW57NGfifsOSje7ZNMTo5uzXb1hlnxk
8wR7/mcVmbM33VwaETaojOmKow8PZkrYXQZxlrad0lJxgUrGpokNJWCl5e5zz+vXeELMcxf0F1gf
eg4hpZGNKwsWkXXBvUoVl+Pht+W+YUyjQ13DqZJg1n21KKpIQ0yJ3vKGF9euuLnpM7xchypCVE9f
vlgb+3bML3fG7EH6RHpbmPz20qupjm/CUjpI1F5qvui/I65B4fbrfnR/hUhwC9Oq7uuQn0UjJaCv
ycpaG6uPLO3zUpFe8+E5V83B/OTKm9yuqAQQmo68yBxQ4Wqfzl1pnO2GIZaUuzGlm/u/XR5OLi+U
s8iDNfPJAc1OiaPpC3sSTkbmAvch9M2Od+W47x5QrV6STBXyHir8LqsuenF4MpLbGeWj4mtPryz/
QdvrGOZP5r5Kw6XBo5a1sna5bWv2SkReRmLhB8GRE8rUdyoI7GVf3A+/I2qAgCtEBKA9g5kYvjge
uTScMDSg4ozFG6PH4OMH3gpuSnGlcKvLcWoFPJ/YVDx37ZQL6AwXJvXf29EwFoZW2m2p/VMbWH4Z
QMc4KyQzq1stF/Jb/N51vJ5s7MQZnfoCgSqOPY6otxYyaj0nDq6U1DaBAgmYKKT0IYNpar7+2FFX
UzEfs544grRBjbH+hqYnq6dWHXqCd6CZVIjDmS8CdPrbpRsPsjKpc6AKyXKyzbwaH5aUS2QPjTjv
OctS0p3XcqjVSN+YFxW3Fuuo7zWbHsNxfxs6G9gKA2YP50qpWkuu3xx8UK+fDbo9bW15MAYVW7iv
vS5GDUKNZsfgioWO3x+3zmQquMeOc662U1LK8dte00cM8k0yFriddaVlrQkNiaLYW/PEl6MbkyXB
QDT2erNSpheg/lNnScp4o05hB/O0ZnnDV9JEW7kHJaLXmrXbakXd/y21g1nyBTRpgcwClHDEz3FB
DY21M826vOUsGyalFLvxAWModFjKcanfK4TvyCPCgZBXrpX/pJC/mZ87SA426TgRi/0MN712f5vo
oHyjmQBaAuHVnCAs8UbcG58x8ZUh4lbAmd9xA7R0r/5DK87xevOu4kxzzbw3O3/RLiVWYVWwizVs
29uX9lHzcZZ6MrLciI/ESOzWwy8di7X3dogWyLZNzE7pNX0lpib1cJh055ByoKpiz1QXczydt0Lh
LIYwcjBdLOGu0Q8CsOygu3ZTfjZBjxk29HHYBF4fAMKzyH2Jqdg9OpNSyOR96xNY48uNfzpLw8l+
43BznlAZo/LvBuKI6gVSQ/lIkX7UvW6NjLO7k0VBu/P2PpaQrkFGhk1M+SSgFpN2coG/39ZaDKCs
VR2S1juVVaSvaC/9k5P15fN2aYmvQzZkxM8YNEjRNtRrPPk3ZbH7Hg9iF2G+/37mTcftB2O3GMJq
7HM7Ivu6cF8pHiLOHit+bFSQvJr1rykcQ7YhdQadyYUgaZcBSjLEFIg8pwldcYdMl1oRB5iuGEOP
tvCG9ThugvNesJGwiFw2IckcNo+ZmtnmnpYK37W6NTxeCRZ1oWCSpDMaBEmqxvmKWvtWpGFmss8M
iF9gde1hud4fNppmtZrLEsFh2Gt5RQYe7O4RZ5/pHGUVyuzKHGygur5ipwLJm+mIM0ckooAaACab
HarAWI5Nr6fh9MdAlzdEP/fCXrclmqYWUjR9RZ525tyTYShAvvDoDQFB9GZAcYdUdId6x2H8rDuJ
FtC9KKGWUtI0dUEhE1FPkQQ403yu/mp7HnOu3yD8kEIxKI9nyikVeo3i/bW/lt6871ya4TmTUE8c
7bJre10woaz8WqQPkkFa/CT3PUvbYe/stDYF2LeTCGCb81XmY5lyLIvSKoYGIV4peD2rcB8/m8Eu
gB5Qox1l8JcpmiJK54z1DsDdd8h3LEMwFoM68PPo88DccBfx5ZJqHfTdSr6Ia06g11Vjexqo13CQ
HFIKCRgkoRxmNkm51m97r3WKb4sZdsNhfeptuuj2aMrJeAJQm+0aK2Qjb6T/KWrjK/DhOKqtl9TW
hx+7cqDR9MpZWl+3noJcE1AyFvsdzdKCsndGIedWyetBzItSTj9P/vhe2PD6setjFCAi/7uhCn/X
VejDjc/x2zW3be7z0ReCcHeif7jsMUN+tI4BO3CQGczkAAy+dzcAC/Q2Ikvf/A5faQfIyiGhWtpT
vyH0naeu9LyJmySIeLWqhSVE1EKT4Gg39IZCrT5rUVjRi7tIg1CJZnCbbvzm13S5DyRkM0AVaEG6
OO+Ple8Rwxx5R7B2lJOYJi4QX13e3J/n4nHzPy3+7k6Vb6cK4uRyrIaI8URb4SkON46yph+JpXr6
Po/VeuZHKy3jX9RQJ+7zWTyM9u4wL3SmQ8W1VSt1Ykj0mV4U4AQYTe5yYDTUhLo0DYJXUldrYz51
ulf9tRlzEAFTPKzwaeKpw3kQ54E9tDauf5mKQjdzq/+fWbmYw2rmkdESp8/qnQpGizYcirZiIoo5
dg/FV61XKEoYYkmW+twueCBXHcOgQSwLr15q+RlcPP/0IQnt5is18MqkuSgKGUW+9Y8kxZBkFJM2
LmL4Q3U4Yd7A+Kp7q3FEDks5aYQuvN0+srXfzPsKB6YYW8xr4jEq+R9gZk5OF6/PuRpOA9J6NTBe
dYo/RGXna4XIgL6+s4yobvkV5ltm9W2mxqVqNJpTp3WpB3SAU/3NX1NJ6zD9ArXRtcCnfhOVd/fu
hciXz6QHi5CLQFDxbOx2Zp+mdACufYMX2cazdeSsdG5mroS4wPC8nSD3AhR2Lz6EwrXvcQGQ4ueW
gzup924+C0Y1zcoS6geZmQIkH7E39Yg2W2rn6/m/fyhOoTfM8FyRZamnftGwq8XZBP/r0W6AeShz
ZWzcigrpj5STfCrOKg3Sk1RM3jEN13xJBIMWrtrxCD2tR1foiR2MZR301+ukK4+JVWXHeVaql8f5
hmUaLWjJ8+capX+5lvOcldvx+JorMX82nfEp5R04RinasxUWbjjZHOyukiw51Cei6PUQqeaaSjVf
Lp3uyr4onuuPy5Hacdr0r9z6yBnGgAJOWB9tNfEtpJCu166ugWXTNYSZk+6efH4zqx1L7oTOVuTY
n8fRWsqsaS1MTIWz9xNz1ZGuly8V4B+/xpYKJl6iT11PgCyFPT0uy74cUS4ldIdVpLyGAzlvv9u1
646f9S4hd9pE20fxoVLs3djh76Gtf4PsIdurKbsGpR2WbnLx/1+Mqv6HSVHjopn+NKpn3VPrBFBB
LmGAHajGh9PAKicVvvYUQ/ZyorWy005MmPvxyCVezJ5XQ6lDoGM1Ao6zZbZAjQ+cQ9KKE6294BbE
aXwePCcEp1B6itNoj9fAWMvy/jzSGgh4f3x1jyWwzaw7ojA9wn02oelfH56VhPPXgYyNAMmtqA+u
pK9Nz1taEkEyP99BDu4USQIsQxtj1dN5Wrx88Ltxoc3GZyUkojgmJEW/eWNg9EmuaXL6bvf6uWKw
rf/bKezv4FJUtuddD+tXkDpTgwyQxOfLoVjdMdLXs+lER1HEOPkG/yYYP0y/Prv+EmddKWn7NJSt
iJhA5GXj60ZtUUMSY66/9bJNbjmCn/r2Tm6tsgNOafH1KvuloUZMLIHmfeH47osdzyqyw6SBiZIV
3XmU7wm9T59q7yR1TNh34FEforMF51Yd7yOL3/DIgOprp9iFOKL4GRTzIV8NKtlC4srkNBJ7MXP/
tM1hJ+l1TtGaLuVYGQwWcu3d9lhvVjPDmcLeI9Pp2mjtbhAkQ8BWWQRjoLjHKUTen9rLGwnOrc6u
jooGhkZ0HwzK4m9y7a+KVYmgIwd/o238kVJJE/Y7XQvjv2148kAKdMDDaIWVd4IWiv7L8BIlwSwX
mZyofhdQO1wIvIdFwDf2yH+ugPqB087gAz4LA7jxHT2jkec9xO9aXldVu/kv1uWDLK4wm+LL81NU
+p2zEnZGsH1QYUHN7GI2VkCsoLb5jyVbFTdsw4C4pWWKtD6yA2xRnUv7GLOZdl98xNxfGqgxRT+S
/aTDRVj2ynXQHUd2GkOyTqSEpF1//GIw+1wS+Kn+hY7j2l9KRG3OskFb9wwpLBLDOQ/287AYTwzE
40SN88qnHsgA+yjCb2j8JNHteg6NlhF8WxIZ2vEkT42Q5LEx36JATxao0QrIGpW99Qi0v2epxLvs
fNVCbLfuFBc8Mg28U/iw/L4dHGtvmqjtfXKQopNM2LeZCgQWykHRnLAJrh6k2wgIl9stYnJ83tcQ
qjrqLNyTts2uI5iP71Id+TROs/zdrWRriP1M3J5lqhkDH+BaRzEEikNLsytrWl4BCRwKKitsXxk/
KWWW34sgfKpwVTWs64G8EcTY+TRpaZ9yUKO1FUeYqBx58gT321lbfTeDUnUMqqqdRg7OEDMPSVZs
CHczTi9SGU3SY4AxAXV6pEMmPy1vDddVpv9oEkC/2BKq7QNQ/+/cic/kg3o0TxAE06UrhLANjYRM
0GknifwxwLHPTkFpR8PM7ER5K/EiHuTGODIyQpkOrY/o+0Z9wB3afzZVWjw8TD2U7Wt6ewZCVWc/
4dMml62sa/IcmimfPpmvAJgrAbN5CMKmA5SLibztXdZn80himsmxjuX969H42Mnn8fZt4AlIAhJX
IZ0ARJlykfozbqjUStrvmMKlXOu84D7ZLnZFsnh6o+s6fGkl5G5bzIPSCqZusWWRJSllRjNFdWeO
RBZIuCrPnFzbtNI43YA0Jfc8YIy9OjCdkicbkrmgwI0wrRh9r4gSRInIgaMUWBbPkljIM5YcHcIE
zoJpMPtqwfugfHN75WTQ26eps7N/ivHtBV6cx9X3RZdPxSS9eZB4YELebMdoVZbLpxzlJ3jFfkwg
nTf3LR5bAua+6EgvW1zzPGTwxo0X/DixroTl5dlWepZYDaKA7C9pESmA/xhP7T8iJUCBzWRgFnAZ
09VkSPdKfRgEF5VZpxfdIKQ3/1O4Iu+EAgLW8oeWZ8m3BO42BfS1FTbr0Zxe/Xm6z+qYIBUXyGMt
8GVvwaoj6PFNlDZVO0oVE/GK2eRp4F5LWcQofZgDVRKdF1KrW4HeZXXv1psv3YAk9YhCPXp4/Z2x
acYlMyjOhyKmbPjFQg1ATGvXTkPsXHyErUtA7X+1cBTwhvtDd+AcQt5YCyYA8SSH3RPpq1UYYR27
+2E5Cp/cpHcwXU1Z794BTCipVUB2/pzOPVueGv88LBDeU7h1+SO/m7tc3FKO4dxitAJdKLqK/fEN
Aq+hWUPc7G7id+jqzN1Y/iR5+Na1yx+eeo+X1ucMsMStmCK2mwjNwMJcyt5VORvXOFbd6GpvXuCs
6OrQG5MFYcxpF0F9NKUa1kQ7XpPnQuM5syxoQroDcQw0nN+eFRGiXqTFIrE/Ozkv/e6sxGEz8ngv
cLXpvnukCaBVh8fkuNvExirhud3FW60R3h1GM3vsVZyrvceGxvF8OFU1EzUi2vihXkDUGRRSepBq
fLrWN0URlQs5tzsECAWarBQ2XfLBfS3Ok//z6Z6uyW4Pr4ZiW0Gtc4M0ePrvMe6JeRFiwin1FTzr
9f2dENT8UeLY5nUyVcvJMbB8jgUZzWZpaVVtY/PdsMGIrdIsJozHhXAZl/KLrntt97TNtvlRwa4C
HeXQdLc93GqIXJp5ADG5rnm00i2vF92poNcOSs2RR/G9ejNIilv7IscJQCZ/YKRnV+6xrQOaHFlu
9Rx6DLyrqAz1gWtlgQQSm/bGJWgHyvmSXR7hiyP+pr8i13t/Cl8OrH+AcMY1r8kNWN1eBn9znjix
Lvv70VGXTKevhqbf+KGdSfdLpkuzFiq9md3JUfOC5VCVPVpPAJ9jJwoPhtodib1ougc0LWx0S1ms
ffl8XnD5K3hHjw7k2W/A2mzpcvAe9okFlo5qpJSBBEcAQWQG53SpnvED4ANE1qBhxzCDlpAVs3Jq
sI7tXHINYYTwoLJDX3+Oo1Af1hP5jiTLRPAmh80pS0yxw24nhN7DK9DhUxRK53xMb62ZdYrHr7us
eXqiz3LOcHxKW+0LR/LS9e+nmLNJji3KubpPnvQcRCDeRY5Ukv50ZjCRQsKIJa+KsnJnhsF2VbfT
F42oaKGPKh1fAx3m0fhSe+CdlrjbXNaJmcbrzw1WNv5y1Zi/jYcuGfAeINTbwhoPhDZWMjzLZCfe
I7lA6AXoU94zGciUnSR1PU+AtsxvupIvff3sYmQvs5RaGgav4St+y8y7/Tx0ydmWCKU1hD0wBSbd
oYeolJ955wpq89zqESmgO/9ZSfjjgq7htkmv8q+qKmr61tK8JKD1D1qCaWmFReS/ryjhzSFlY7Zr
McNRYmxkzao+uqzPe/7ktHkmCP699jYJSql0IEdL0NXYNBztWW4PibSsL+1sV3dkK4N6iBJBzT66
B9SHE3R9SYqPzbTQLYrX/rokQGTPI6/N2R46woKQQEzzgsc2QWbhqr38TETSTB4d4t7K0A7qZ8me
2TOF5UrHGzvj3+nHIgoTBHftyM6S1QfR4pdwcbCzihym4h0YofYuLI2/zFJqazJiYjrOmbVCM1dd
vfQ7tAEBuAGYqkG6F+lsKLRZssalefNZgOzA+Wg1c2RtAmBNKJgX8NRWM9YRmitCZf1Ug0WSylWh
QAF80aE7wUTp0P/lwbLD0UrKLXUP60VGtBvk3mUDh8goF2ly5KCyy4K53nI7yloxpMGiM7KTijLR
s0DTAWo7r5Bi1cMtBWJeAeaLZAM1Kn20jgyXg3rY4fNtaoKyQmhKUhQo3V45jwFPtcO4mUBDPHOv
CsI8R0U/Y9z4qu/tVTT2BVKDiFiOVzk/Ga4X1oREXYF6XnsfI2+3AnsS0stA+Fq61FFhLuatUn2z
08I8fTgf0hkLT2rJzh1g9FecXN4wBIizHR0miXn007Hxr71Ag/ckau+xo0FGAhui2rAhn+svhVqI
xd0QVrGJDmfoMBkd/I1GKVdbIutTVFivHP1Pm6NkpKISZfYRL6rXGHijuUOAT3s965BwNc2UtRDW
LaLMR+wZ7h6gpuU6kBbwiaGlKIklBtHsyGzaz4kyiiqTlYOwWEiSaeex+xLckLqfnLwjMPkw1q1C
xAFg1swlxpQCieUhzh2+4i4f5KqG9g3Ax/c/USFG04kgqsXxCXFAKx4ShH9KAgWHyfZKTvJGMQxK
GQ7YWaCE+7hpj0KYO2a2zs6SeTfW3QnQ7z8htF9MUdXx1Rogfpv/9hdqY8OwRTEI40QA/eWnUKZq
sHVbK0OBkXPwZGBPN/Iv0xFzGz+QpWmkqDPmfpp+Ywa6h2r4E7rU26EDm7NuOUziJhIYk94FARa5
JCi3wOytAmehOSOFVAMbfnkysR2oqh8o77RQV0udHAiUTCySsHD9JEC8mX4BHSsTDnGJ/nV2bQXK
TBaPR6bbHhNB68GF7zwiFuy0Vjn99LhayNwsQhVl1wQPPAgzISOckT6l39GMYoPWBG9QolpWNQpG
I6O51LB2EdKnnvg4uMiozOfU/oTbKJu3y17zgWXffUxwY6dlR+msFtug94TzVmiJQkwS8TWyH5to
OtjpgQ9kTFYyHk7sUgOprcfBqwOCzhZPUeit8lYXype/urW5gn/RFIxLmZH/uD/CQFa1vmOeIrAg
0j2iWIvlFRk6npfVdswAO/nW8eB0wfh5IIv3QQL76bOeJtMxmyLW1fXfMgFF1kt7u9ukcpikQX9d
EC9ApFVQLDfIMhjxg7YXw+zzGa+TPt4qnIU7UNkuYGni+ZvaPfVK/xvlhKR4Fuj9fIRfoXlLnx1V
68via/XESyT+Ti6buiftMJx3iERhn9XFCw66C4wvWiI7nXPim4TcljKsDiwv4yB7UfcoXJ1HWzIq
QIvsf6XsioUEXT1e0/OdHcq65rVJqoS19oDuCK/PhFOOyfnHHuwtzMg+/UNH+ljDnAgtjCeUpCj5
+6mTZjSAJ1KF5BwFw+ZFu2wUrN/VHxeNsT9MF3Qj8cw24jLQ926y0OFvBJd4E0prbgOR/M/8i9Gm
hUaD9cwieTb0XeJMxiivqulOupwTzxmqSL/Niy2+Gcensurr/dt8AClUHpGciVTMhJyzWe1LNSDR
rldzWH6FPQCXQ+vAe5ekfam492WJeC32RI0V9gCVVJuMh+LjfXSO0OIWxejIgF+FeY43QrMWN2W4
r9SRkPBQOTdX7nO5jF5YStkHkF8C9BQzeEGyMk8UCtl3ryXZPsAurl7yISgHt+/UyKjCzNs48Se4
7rUf4KUp3o6lpXKKwpBvkIdJ7NpbkNJc+/TzpDR17Ke4d2+ujz8VsfgQ8Vt8Nm7lzDfRT3tyrnNu
5QELk1LhMsR5+IljyFZWaAbc5qpLu6BI7LyOHYnpileMwBoUf4tvNSJFDjo0EzJiu5mQXNZQd/SZ
6Hxw697fV8Bhy/hD/wUZHbKqEFa3GK8pfHMEFJuZhz1UwsPvlE4cU6SSYgTRa7/g+D719ihxXur1
V4+NyQY7WIXBqAkeeSpOA6AoT9KXP8GD2XsmuyPXUhk85E/BaBbQXLvOfna8aK9TkC00yDJB3oD+
ggpMoB0F+t2gZNN1ZZPGDSHLlld74BULgeAkFbz4F1P9wDncdZrP3RUgpun0ygLlBy0r+tHO4Fn6
RSetEZ51pF6dBQJSOYXMSy0IfFL2WLOFR+sMW7oFtvzz8Q0JwvMARit0h3k6p4zf0G7GjkDCwY0z
9p+ve8Q7lE9o24ggYSsAk82nbX/di7sAv8PjgKnFr+i9oqU239GPiiUEhNmp6Y62S+yCGxMOZOLW
0WhFFenvh2JEPEc0MxHlQEl5tenQoC2JR/N1cKbM/uVxCHxsynjQonBBGtv/fYVVnL+utExWSfIi
eHTZzO/FqFbq7a+pBIJunsOng8g/qp2Oz40Dkz8XPiKA3RUc1OJbdEQl32KLjFw1EYLeMeuSdcL7
GAe1RrxICCqs21GRYcBI4pLquTpQ+VTPJlXN5GEvoP1ptZDqGOqPQxYBWY4xnC+R8aY8lDzewrtR
+ErmXam3t+7HED+YOsVmF64ltIK95na0pf8yTjWILWxa5RDia7idtrVayt4GZrU2mcp61LrhpsmU
ooat4lo1L5vjY5bmTYBs6pJGkNKVBkbuBhDXkCD+7J+bz1u4HIq9JaGHB2HXPgf0XPQZXZmb1fNL
tvETm/+PIJKn2ICm0PJCoZsbXZat94W/UE2ojcG7wvpF8HWVaTNkRi2sdzloTfWJ3cxWPEYwBAke
1lfs9r4eHtiQ71P08y/I2IqX0yIUHRG6PlPHEm7+N+fdwh2KKf0NJTDa1PFeeFMytulb6exd0pgz
5oVPtmf/OZ7HuEUBRHt+zvvu5rguNTj/n7glPMI4haSoEmLWe7kRdchu41TgiZVXOERSIaKoXrS8
g2HjA4VKEG0SxpZ6fgIEe+ITPMDoe4akPwkBiG1gJKe6i9elRO2hBW3MAREdgv+Fg6xAQsZoblln
iXwBhWXWmCART017clGHmLdNvHJh3y6t7mYQyAazqdbhl4/QS9Tpfh2oLmhKkSHNPdj3guQZ0Keh
iYLJI3L+RaHN1tT+pHtKV3Gw7T+uDYTkv4EGrWgo6Lp1eddGgbE6xOiCCkc4LUOrljGtU74avuZI
f7VqY0wUoYgHCLitJB4t+QS6nOK4JVGK+l7BRoDlUh/T+fdpNO7CHRVOfizf2aYMyWResGZTgsvc
+DEUtoTItta5jiKBZWPuYOSPpirjOGUwUoFeKUUI4rB0vjMc9egcFsaCXDv2DtnI+t8k7w5ntvC5
ksnbDF+Bqsu40YiYkklz4ytwNkxDDHTwFQV7igNui/a74JNOFbccdhn0co4MaGVUx8N7l/UwjqjH
ygfzC+7nhuqas6uFYYkWhA7kDByVqN01RLPtCLDjC72uefSLT+8HE49aNKwahQ2B4dlZaGXWKGXP
8aYXERjBkdT7NB8Ruz21XMTz6wUMoEWsZ6ghEtTJ9ws3QEe7UTH3DTAkUIrZd70xF03laaPe/iAt
Lzofh9/XRLK83gxX7Ep4x9mb3KVVbGrWFfuZR82SY/7wJDaxmBcHeE1ilzRC1CVUdTewZMVeqM72
MKhDkocXKrtChZ/q2wBTqUG6vE5ID3Wm6Lt7w0ggsPdgH3drdPjhkJPhEP2r6YY0DYO6YrTSymIO
OOFahNQuBCZKxHPpXyHE8rr2967ABa0auvGbLIfX2wcRe1JkRctIe8dAZUI1ELiyLeTC/V+47yFS
HMBoW0Zv/DOXXnTxEQT9kWBjzF3PPK+GH6Kr5RA0Rd8HckgYmTsL5FbdPlGD2+HUWW0NrHpOThHR
1VKpCRdcVNK83uQSdIKiAbhn2iPSSuM/PHE/u6T5r5a0MGcudyDCgW47YNm30iCNgm8d/Tz5R0kI
rK7fCmzOycpABZDjeFofMbSbzDzG64AOykCzqjPqtJ1c7cJ1EkjU2O8rRm29msMxIyGFwpd98Xvj
deuHwUlSJhbtTZKi6Ox3JvL1IwCNpj7xV7tKTCay47sKO6JcEowodP2RgIUVCb0euX/QaRWhwEx3
4u63RpXy82SfVrFugNMVYBAxLoPEYN1v62+ln5OPoIxa5Xa2jdOVF+q4v1TbFmENjcbJp+NzhGom
rZnBGbRtGMs689glfrl/gQCtwpTw6UamBIcSLP/MAt+emZfA1Agm8mQZE0B+JH24aaHRqxErlAKl
PCf/A47ycXqahKgnG5FftX8f43uMImQ2onn8EeL/3k+qKXU2dpMhzCSUg4AYFbOIi6XrVMOLoVOe
EDpHSAf9oOD6py8X0hzOV7AC+54w78jGuSXb0WozxFgfhUO+GXGvgzoe5mmAfLdQBhm86VNquqWX
gvRo34mdOCOPHtMGV5T+m5xzLNa83GkIrrvrOZVHiRwqiKS/qfGhmPTcykQa1NsI45Il+ntjoOZh
xXfZPGFx9KMmCOYzLfGyxEnaHUCUbHEb1qREvyAiB0VVAsYlkKe3G8N8V2vdNG12b42d7VXUch23
ZHfaimPsNGBiAEHAKA0NQw64Rz+0mNNjdPw0Tppi5EViM0IdbAzQ8BZhC+tfqMTXFeyGgAjJvNs5
ajUHFHlpsnrKCbN+Pq/iHBp1fGAi7izSs9BhB79y9HBIp26E9LrX2WA6d8JCfIkTZwRIb6zux2XJ
MJKfBtsN5xtg8Jln6tENNZeyF2Z4KKl37ICPsyMQ5OPa5QI/+RaiF1Vrt8Rac95jXkXKvmysgm06
c2E/Z5U8SrJd6dQRevGSTnNbBGBdTTiikExuvPPX+Tn8Q7uZ4cFR3LZbwAnFch4i5RpxmwJI+Dy1
2UC7UYMOWCW6bshOwd/wJ12uZEob3QzOYkJnUz3STrhfu8ams75vAqWfd3J5rVKM/O39x3dX/Ct9
9yCJ3f/IbfNgimYKO3b5zGVx6w/ortVVHFEcdReQ8/qwXnRKPqW23I7jTe9X8RDrQklxuNEMhJFH
COSLjCMkl5WMg1YC98meO1dmwT/ojWwqR797IEbUzI5QTpLsq68KNl/vqEIHkn8cfir+xwT9QYII
XVBmwaXGt9gk55ws3LtizvCVr6ShDtZIF7iPygsVMdnidFUiKrE+Pkh6ymNYSGg8hn5G83/UqmsA
/nINcBSg6g8ev28WqIHoGu3KBAFpmYzj0d1Qhz6eEbvZer1mFp22s9QMcjYVFWdQUecMolHzbBdu
eNE89s4Bad11pWxMJoY3KbzsG/qYK6IlKY5dGini/JuRJnxxJL2B196Jftv7rLytCOioSiwgJtcP
OUXTX2r93tVUMPeZzOO4kVJ9beE9PLlkPul1/QWYzfGK/PWgl8fewAwi8sdIGZcPeSza6nwy/fxh
tqS/WkplFSo+JqWKl6UMVavG4nWf1XbjABVm7m46qDnzicKhapT3K+MgTwr+B8cLlMujgL/xlqkT
n0xdPdZPGPLge6357ZCC9Dq4bUj0YXjfjnneFIvOf+5vefWni8nTfx+AzczWHuw2+Fg/Sm5R8DSZ
kM/B+Md8d8RSqHeZNUV1VYyACO2hZHPAl8ZLwlx7dvRe8K8w58eEKoEDWILMYejbgKxA1YwTKdjy
RT0pDyZpRHfZjw1Hr1tysX+m1SN03YMh6UIek+sZB9d+1dclVM3Uk1Siikf8MhJ1QaK/nu9kowKZ
M8IivT2JAyUefsV4mH05nKCIqP39a/jVURgW7uLeE4TC1vepvD0D+ptiaPnjt88Rjn/fws7UUBYv
WvFepUt56u9GQ3kBnEP/n5PzFCsjaaDRinWwELhD+fnvmGL3dm0c5+9bsnSCQquFyb3FW6dr6dZ6
P/6qsk6W9fFDO0lx3tGIz5rZcdoWOgTO71/reJB1pYkL5Z9+VsSB4mEfQswtiJHInHX1lkABtBDA
jNilkO8Pg9zS8s5nrJMbEtrTIvjRSbjxWjpLI62x0rCdR9ZMdiSc1vhTJpAn28UM+8TMlCIrFesa
Xox3t694ngGZxd/jp6z5yU/GJTmNNqUPpdr+in5hOKwAVOZ0H94l1wS0dUbDSC7iMXd37MRYkrc4
FLl0B6NkAxQFlQf4u9DL3vl2iW39a0qM7nqGqU1D1800AhXUE9MCw0OV89DJYuzYy2QRzbwq+pU/
gkY8L2HZGUewhpBUgOaI2Ab/XjZpiE6ZFjQo+YyOWQi+wIGLbmZPEHWekvLxQUqsmU2BVjywbGG5
3B0FT281s20QL5dj1siuy0qmO/mDtMWJo33SUf48aXW59ukJSlyyqN/NB74E5z5UQz9OcnI2hjVC
SWeU8J5ZSIfzQWeRnbFAlwUFN151ltpCTsMou0DrNnsE8GPy4zmVROsHmU3LKdbj0SPdtXdmq1ja
WWR8zvILIQNhzOxtV30wLHdwelMzF8oTRPzJ02/dSZPQuqMXAfVU5OwKrcVwP1KREEU+uBO/dDP4
d1KWqWaAvfRMfCYBvrHXKWyhF1bfU1FEYVOillG5Bytw7gLTu4a6ImZ1El8BM52vrP+DpIjW3TD6
BwfQ713Yccy9vqgO2SZF2/2miUp0Fw6lGHRhMrZjyM4IW7t662J2IRWAqqtVijYeFM0njoS8KMpk
pv2yV8pNWnlu26p+EIhhBW679CXAJlvOpErIGNoqeKcAkGhZmdFRRpdX0wnwlAl4QnYWM11W1D/4
c7VqZfSj50N1FknrO2xRfyU+9n16D1z3OP0bwIzAwtxKLkF49JDFQrKoHZlkqfdwKeBN3M9+Hanv
vN7ca+w/53D+sIErfSSYoEUQbjHJdopKVkt5+/HqDp/Cgm93tmxP9u+30ZDcLMa3zXbuLeqlTmvT
EzZlcvF58UwRFPXjS1QBIn+wViHtjZ4MbNscVzAuKbbV++PGvhqdrR/Qj7MbyyZGukMxI3yn0FCm
XBALKbHUAfdTylGfXjcDw3wOOQxB1rbswVJvjA1T+PX8bUpDmLTRv6IKlVt6UkIHNtXMKL6Mh6RI
DxVzCEdOdz6qUq+6eSx9ShieWmTomNCR/Q+A6w6Tg8O56aE1s5dOw6I/08srrE+Ju20vY/bEl6sr
D2AzEsuuemNssmEMV4IEgDe3YqPfq4c9pRbRJUghCrF1Y8oXipRILynVRGMdkF841jKl5gxMLrse
MR3z6G0BKZElB97J4+XHJDVrOgMA8/5aj2swobMVlC77c0TvVY4FfbKm67u6DMSDGXPUnE/ywoJc
+85oUO0BEgHhwOA+xkpSzpiIpQZpyBruf89ZFaaO/PNf9+3TM5CnCfM0jLxYpwrgCvd9fbyb4kKS
GOYXcEqLBjyt/C0y6MIYa+043xHUdJPEER2HejfMPhBDmCHSlGecHGdGE2oTOREFMH2x8lpf4Zjc
JTWlW18QMG08HUzfOZKuVvXuzNylCihkiusul+R4mKAgoE2Ahhivta2N91rGlcClJaeY7e9eyFZf
e4yZIiNrE14e8yUTOH1Km9GeBoRdUcDls/jGFVeipGij5ytzXl9nzLlKr8U5yEsAoIcYdLzKvPPx
75GnVVZBfzauR40tGCACm8Jt57Js4MYRZjqmlSseXm5ugiRErXHE+IwxVsMBGvp0vphrVVi54Ob/
7Y6cvCBRrbjG4jjNo1YkzLlgJfyPfQ7Z9eWpzDL7wIHuGKS+DO3SE9+sGgw0EvoKYjcpLkciIFFJ
ZxFkFrfQrEamLSch14PH6IVGOUjeDWujeJ4p+oNNbbHByNky2n1V1oMZNbDLSN8a07FlBv/d4Spm
9U20Kc3wbPa6JGbtpairS+79zreSzPVPq0134F/9s6oBtsPoCZXIia5bH55m+TaBs1qx9SrRijOx
Ovn8J+DDLsuoe04Pclo3+AVO7WAngoBPyd/s7HMSq1NeDAmtyDzHYRPapVMlin3kczNTmO5aekXi
ePJz6LVH40N5hnSXRNOej//f/nhoUkbzXtI1A33Bd3wsPIgrZyGA81ZmeUD76/s+vZNm5c85/Z/v
EvwjlN2yU3j/rNx3xnrGgE2xgqHsWw5PUdB5MEGPzSAsrIzarUc7x6iDtCAB5fwQTz6W9nPJVpcU
WbWxn1nNMb4swKpjI+g2H5PperDHNGiRqqUycHi1PDpxji1Or7VJ00btoysevERcjo5W1Mips2+0
f3B4q6RbOjvGmzKa7WNAQBAbJ4ypBv54usxiViM2NDrJ/mBo4lTyRV7B60fc6XeANFxdKTMXj6iO
eesrRVJ6KYRhBvn8DKJIwg5s1FnpfJ4Rm88zPmZnqZ0m8sdp7FbUHrQqt0iMN6JkAxWevtLCuRkV
cBzNSGJDeqEXf4v6Qnw6WRl+rqXSfoTopgutKgpxZ2+tieGBBAD4E6lueGeTDatqxXlGElRl7C75
SplMxxE8f2gx6t1gWdAaHHXG/6G8sURkAKBMtkKOmLvCYdBaWeNYdB1Nk4tcZ0Z0uNiGpgEkNTxG
vK6YgnVlaMdI/oYAHH/6nmVRBMNa2/jtPZuvuZ12jMlIeROewocVa8AOL9bu14YAKV2t+sBNsFY0
a3tFDLaw4eD+ALgjpaGrUVsaoHgsTf1kummg9Yt6TKk5cBgsolvkXEGgJoCP98UqYcVJUrwBoNWe
2kCtND4Om6ef/8LfMJZfKe9uVDm9uJ983cGy+Gte+2QvTz2Cmym8wjmT1WYk6Gox/nJMWZORdlUF
LsMwBMP4CoG5Xon3AqjjWLa6WZSzO7UnghQpjIQsOPRPBFCdYNLQyJTm9W7plsOiQkQZ2ZP0Er6Z
Qjj8bUpsTdei+Bn2bGanMws6wwHb+hDNYQYTN238zgeA8eXbR4nj7Q9u9goCcuMIn0Q+GIGXg6OJ
LJDMnWBGobZaI9JnMsgbXSa7ktNjvxsHLAQISsWaLlA1zLJ2uTv9xBk0SixKnQnnZMoOOuoLgv2V
R2ep5qmNWnhsE9GQ2nRExUbK4kM2T78r9SCjgZxYNPi6TnE/Iuc482SImxJv+Fc+HSyUfPXxhyDB
9FKqJldImVKZijnXHamaDWvnnfu4LPA9+l46ThngEcxBgayoZkYFptUCurrD0ALBFtVKDuUrw2FC
TZ1lvcYDpI01R3Ono1b+DVI5xLFvDBxMBlwM+ep2ccWq+nLd58g60IKYLQvfBIiCxw7NJ4+To3uk
JuLQUVli0/v6gSxEh8FQpsfIX938dVocZJxBZtNUzL527V0T5txOJdybAVeN2n9R9WlElIVFxewm
8AKZ9jVMMo7VZ5xIwdcrEjkuguMHd4wtqfKvas5QMB2R8MJ1+NJ45O2e4hAhJnQGnLoaLMr3JQXO
sQVIlmI3eyGCs2pHUSRoR2oidEqEOM8vGAnDMpMvU7lQfUmwML+uhFLtYaWA95xLy2p3CzqcFmN5
CBaddbBrVjcPkpzcom2NlW2XHTGSiKcppMQjFBsi2tD6QXcUUyNBylAY+IKOh7FzJZ6qJQo5dpak
TiI4g7OldS+nd+O8yCND4VaxxR73ObVI9k+f3CrpTWbuGg3xoh137prOl5AahN0fwWYn1U+MjOJr
Jk8jBpbnvIDyueKHcvABARi/KuKm2KZ3pO2JTwrEPR3LFwBJu19pQSh8+/9HH69GaYQyIsrz0+6K
QZvob8EayC+f0Rgq9GIrI33Tnj9dV4zxIoZP0wBOvA0k0PqCDgH2v9pUTF0yS7lQ+ZMh2CN9iT4a
J+ban+V69AnljZzAuS5tbZRGxV2fiNaAct9y1QNcB4k56PhzCfKyi1uQiHEOfiRTPMFNOQkbZgcS
8Bq/8BzrDkbvaxOxSC7JHplcSAJFbTrCaSu74s/32MUb1jh5D8F4bAZlt6zne5gg8+ir4U3CVg52
XiHN0Cvg6fyXRKoGUIvNXKRPQWDuoS/Iu+Sf8hh9nVOz7eRAMQcmaKvB45Fxbzo7XYJFLJnXHhfz
yMgUgj6D80wmbHW3GngtMZzavlVMmmoeI4a9amzE9fa5rcXI8QRfsLSffc4eepR4g1Vtw3fvsVZg
XxhaVaLBBhIWxiz7oj9ccnjW2QM5rvQWERcE0c8WyBjQ9yF/EXOaROf7TGsig1LpKwwgAZLo8v9x
fjAMtCE2K6u4fPW1UMQzyepEBNrT5edlni7yzNgavzn9qb7/6wyQcQRySnUsPT0b1hcZ6CpZFxv3
gJHwhpZuE40a0Yeo8paKovqTD8b7ecwPAEHFbUAKV1sYx1DjQEfbsDC4wHZa/+tOj5bq+Za5hHRL
8WVEtG74icX0vkQZOyJjYq8gTtm9DlVoFjOVSGuqMpfP2VuBhc3FAFB5+ifcLuNQrerLFSNsMghR
dGTIU7Aa0VAxh+52j3o9cpkJSbXiiUqxgQZjNSZ0L2+ND4cscAfT/XWOKktn5cjG8SUs7oZrX/Hd
2fTzhD32dEm29/rRFM4puQcCOisFMNSU0cSLYpF7RdPDEm0taMhq4hCfeyU2tLamli3iQWiF/VV6
BMZfTti1/h5oKP36tFkSdP0GgW/il6t/+Nb3eaTZKLjA9O4OLeIMRtxBJAx1p5xRmJN9fGSZ6LcN
AVf87RA4t6cW5XsttofRLcgryxLtLyz3WEN4q1+JznGRc/mzi8rJYzeCdGeT5r8d1n2QuYY6jDTV
5B1JRB1LARCfwTteVneZ/LPFg3tzW2ThkQgr4k8/JKB/UE5dIo60kSsP1x5ahn9ptYsAjlxArnG5
xsKPMBYzXm4UoJMnL6LmaRle1cAAK8NHPl0J9s2vODfbrhgt2FWqUnkDkeFvKSO5gmd0rryvmIZi
u1a4bI7RuxSUxCBfikJsWK50y32LRNJzJI3Fv2ZlP8iLxE/o8gNW0N2mZmxmB1VZ0qp/BSwF3qhz
Anx5zhZuPtjIzGQdgnYQPJZIalwdGz8R+vBaVNvM46MoKrdRpCfPU17jcSqA667xHKwTh/+7kcAf
1jYkxgRBYLhWzAaJY/FThvF06sxvGv21DVPXS8/Tuy5U7ysF5abcloEP0I7IArTSX0kg7L3eVawz
G217m7bVJXPfOn3TU1YrXykwDa8Fw+OnuD7emOcXrDCWoi3V1+CuSZcdJCDkMSacW63Lt5g3ObvZ
6JDly9DRv9e9+QAU8p1zNAfI5qgmqnGCfND0l8Z0V9f9OVX5hUf+WaIBXK66k5VSPNTuHxcevFW+
lHrKk5rM3p5Y4UCeMxtlhjgiuJlvGvBS8txgDVV5ap2kB6HDd4uefL2thQBJdLMjAPvRq0f134Eo
p3O6TQMFr50jQd6miRJypyReX+3kz/UVfZ0+iu2Bgqq+bfVBgAnkOD8Jw2qrkwtp5LMWVBXtfIWb
dHukVaVa87ZRW1wSuNPBXRirLs8qwUlHcxPpd91TMU8bIkYLtI0UGUS2W7zZQ0ACqeM8I+7j/kN7
KLX4prlUEha73En4MZ3ux8vBxuqI7FMVaQQbQy+Op1NvInCfxwTnmygm28dFlcfOLW6WH5kdGqS5
9sFGGgBI3fEWOkQGFLaEfqe5GE/BRJHJM4ZsBHuH3uX6WoDPHy/mCXLHfiqbovovFVuzB9t2uX5x
FbyZ4WADjTHldt6+5Crbpm1Sa5PWdabyH3Z1mg8yeXtrTcKLrybjSFTgp3S1RPk+8MPSD+YFh/aN
/ucQMguTnpq/L8+NLHrvTZLu5lazP7HHxnpdo8p2RcCr82iE8VHCXEE/jifl7efryQbFo/vmAckU
wzU7jJFBW5FNUxY9DcAwjiNP+uLMXDj7gPWrwXoZgXHrtE/fx4a1o8cYvsUhYFVLjonTHY2c2cMF
efexQmepXm161rryqR241gIwKJGPsfeWqBR3tegawSvxqxk8vOm1tZ85rM42ziN0rALi/YywLOMg
iVWQNJ/kxIgUJAICncMs33wVtJ7wnsAr2uHxaUibLXaA1X0eiAfhJWe9Hx3Y6AHGQ6QoRiHyOWOp
Dwx9OndKIXUf8eeHffxzECSWCvs5h8guGDUKsll2pUQq51RWrHDPwvfD9tfPRcRZfV+IrLFea4e+
cVziR9fJq7fznVcOf4wmKKLt77NmBNB1jHBXaaYhDycmLQ5YkJxAJs6xQl+eyR4LZYkujB92TwVX
mCYK/aOQ3zHw0WcI8ISWPdYocX8UA6jvkEVCh2ljso6ZWiYkme2agzDmO60xIPM62hXae3nb+zRL
iF7VuqcQ8SMrjH0FT2MMWdRAf7HRtfTjNXcpnguwTeAkhhKAkTHNHl0guEd81noKlkgD5ZEsiOf2
VXoZkVvDNMaq4IFw+bFNbuB75N3EW4Uhfrt9bygSIPhAYMYeN5oXq9prRBHUXgWF1dBz5r5yDHoN
xA9gX3i26mnXsF4sB1B3BhUqxX5xc/yyrDaa8w9bUDfVW4pRmSQvA+l3gGfnFfQPCMjWy30rfcry
LuTNuSpHy7E1yIAvK2Ho9CzHCHPBEbXmJ9ykFS8SVF8wMp8JaBliIqbtpXnzbieWqZ9rtiUXd2Ey
Ise5jzIlAI5z+86D9AJkjITh3w/S/g9zZpsUjWolt+LuORHw42GW042cd4JwpB87pZg3d3r6B2Jg
AzV7dwg0JrPIY8RYPyR0umSLZo0LkuBlXopuGE2n9BFQi8pNI67O+5eUPUzNOBKPnMPjWiPIVQpx
pHbftq3cpgIar0ggoa+fqnDDSgxLCvJ4DkpFlKoav3ozEezrgPjZkYv3I2c/BskXhrdw6SFQQWpL
sCHkg5KYMVfnJuqQG4hMaOo4BEZofiSJiHEtmLJqmReEoeurZG7TF54ko8i/ZH44iJKfjQYXbyGf
YZK5tLDFHHP2ZQc+v9iXyY4nBRcfgqzURR8+IPWc/wqtzKUW/700cDrctRgW3DE8mjn3XkAKunF7
K8pQ0/9S5yV/zwkxLpe7IE/+lnfg+g/JJGs8Ux3EKfHNnCWriwR3MLd3oKBaR50ZT+GR3mivyJaP
JEzyWH3lwtK3dI8LCoDOE9gmsvllKq1ZksAo2PnDSpOP0HZpVZaaVhWV1GboAbm4wbzZiZLmp3cS
wBU8oPZj57kyP5boQP/ZJCt97QVJyS7w0BmpoRS3AI15pW5zlBEid06TLXwq9JQWZWPE7HfMtYDK
wKE/4P40uPdKGqMbRA9emRMZLyD/Bwlt/cUOsatJc8N2QuuRpIGuQFJ+eddBV3J42xdK1viLzaIO
3QYaAepNcPHOzOdX8HmWThuUq68Sv//DbttkvyoacXumuP2VgJicmV0l8AGGSz+TJkxiK83ryLLl
ln9jUTdNeGm2Y8hZ6vA2zUTsYsciIEEa8O2jAC6RZ7wJlQPTEHmu4o+xBgHpTc06mAdrxZapCItF
VJ9vDHCRR5yNZacq4Ys8YYMK6zHEcEFunMBvFNwvM31gpcL05nTW0XRGe//Rye8edUlwDmmRWb9a
JUdcqlijSkSFhuTmvm4ug79YAvyh9NNKwWJ5xA6pe9Wm5RDiiRjVqR0XUL5es51VdV7l2c0VqFo5
K1r5gx6qfv8XmuqMI28CsVzFNHOcZ5dQzj9Lyh0DwTo2UtWdwd8cYa7ZF1ZbFPQjsYfxkUXpwzha
tEtwFS1X25dUoaKIVk6bMy5awOLGZOLCb6p78cJELDQK2wx4yRpq4FZB5dEq5xnIlnAoIk6pK8Rc
64IHZpcf713wnNbkQvmOQpmHWdjuk0b+4dqi2ZwvdsBMmVnsSRXxuxjPFLoJsjVLjUKUtf3RZklF
tvmlIafXHTFvuKPtKPMIc7Z9/hauPbE4VixsnNRZpZdbT4i01QFLJbtF7BUHXpuMQnqljGo/mQJW
4tNSLvCwBA1biLQq8Qz9NrMwG+69jrqRE4BSdLLXTpVJsjVp9k8fd8JXDkgWOLPVDIHQL+9Xn8D9
IDyfoAu7zjvwdOjQMg/Gwya/ge53YbTL5GqOVEixK1V0hcIq8bZtlrz1HifQjx5kDT/whW7VSsHQ
96gmiyBC058T68vW9EMaOvAIFojN7j2la6XVzRCmb35Rum9BY+rszxZoeBBojVRmQdaaCK3VS9dY
L86NzhysZntM+dGozAACmBb4cyLfW7VFUQoC3+dU0Zi+lcPGevVApT6sBZLNQY7nVpTfwqv+qzEt
PtEfAJ6ZbZ77GqgIrgA0BaepwYg2NIa04topBAOVsLqtVJBMu14Ag1LLYUnoV+KT+SiHnRBSLDrK
WdwgU9zHNwFoWOhCKLXBG/8A+fY/TGT2mM1dahJKPHExa8mh8cPbg/NAlv2bQE4Mos/gzcLhu18p
8nS4Vc8nxvIkMHfrTVdL/BI+xuVbc9tT1kXpHqezbKGfPvubaCAYES9JJd5EpGWkOvx8OvvdQJMP
6aYlcyxTVGjKwRlIsdK4aS9NAE8AftjnP8vdSYWJSULU2YP2sxM0okmjAkCx5epp1V9KmXSgzwlp
e+OmBkMNZNokxSGoaIEnpWlcM6p2JX9St9Hovmgx1ItCdsovnMKsnZ3i8h+SuBY5AYbuk425E57Q
wWqNyX2euJuWOB2Or7pPcuPGJlLTVs30XY53a/mWg9nlAhIZKJmMLaPrKoyLUiPWYt3c/YbAz8PW
5Q5qz7SRg38+UoNWXvfxeiUWwpNJxLOchI/kr1jUQkTT/2c2vtGqcsgIRN/Z84Bp9sWzMZ/J4+Nn
IqTblP59c6N4pdv1McKSjMtvXxEpCxI9xBTVll28uNeWScZKoT16luoASPeS4BrzE9mc8leo0un/
RyRkY45vETElwJxrTQH0YNrEmVcLMc7LMoAgb/oEi8OFFitMOAtHnKxw5PC8s2iuPbhhuMYOJ+yJ
+h3HDSgUD4dGPvxIGrK68hmdBqdU/7bEBvLtVx80vMqwyHzC0a9RoLPLuOzdSuALI3Sdj2roslrW
B0/6WpGyjBwmEZw1f6aCwqw3iqNhjTVWAOFOQPh3Vq55Vr5kKnQSOqfWAWcjr5m5M4pbEdyJ76Si
zqz3DZb1xNMgqzvs3Q+L+QKGq5+AhFnRljpIW94b7SWYFiWrGGQPzdlHDQB3JWd/M0vKnWDM7TdN
grw+rDTwuHTvBQNUsFnnc5nLxDMAx9dsFRcu3Yqsj3M6NCu0Qnk1scNISmqBkPvZByzd/gHGOrgJ
asJFJ+ZHrPMtzKUwiVkLqiCgmL8xMOyXTlAOiwHk4kIU0JwDP7AC1ZfmrPqhvmma/27FSvk7raVR
655clq0cX5P0bxJ2Uj0EbcFGAiRMgWULdL4ZYE6C0xCdu7luA3ySkS8sThyR/aIgvOm6M42B6qnJ
+7KcCHfLudNu3ndxXekn9VEavYeMFPPWEaXRgML/uHetjyRwZPoatFr3ZqtRMb0FZKiDxGfo8t98
fWrs4fCKOi1R0dfbjyywMPekXMir88G1TmhsuM5nF9p/0nLGFjWLPPfwjIV4nIB14nLcIjLkED4B
fO35C9TV/8MQopBh5zy7IDyHNFFtDA58sKo7RbAvcABhj3431XI6hzNE2SfJ4+EoBpxy2C/sCsj/
exFhyzaJZeVwMNB8Ekybopm8P+DZS+vZPwRhJ9HLykg4cGljUEerBHBcLNPXFCr1ZkciA+DvzY4e
wVBdh7sp+1CXx6la6ifoMXzhz9zW+cV6gPdKORINEFe7KKjGOvyFFwB6AJfzCGPaeXmvYZt/qRFJ
J11Q9Xz4YwB5iP6BqJwY1K/P3eEOzhh/PdAJHRpPSAoPS3fx3WH3Le0PQE+bqBVerl8JeOyFOCEC
nxjGleHmzfjd12PVxjUj4rvDY7fsMce3RZm8zT7KY9fE4xUw4PKlLu4jT4lUYncdGZJUkYd7tFAs
IHb3w+KdatpIBWirYGDc6DjffwLEkJS1BuLdc1aRFlI2WiX8enfQxmnaUbbRB86mlp6eJOO6MmND
IiYn871cERRNr9y85OefYfcXX1eUTbQ0W69zdTqukg4w9ZVxUkRRWpWL3wfPYLh959yegmtCqkb/
VpF/9zQ1AA9NVifMi5jm3jJXC5X2tkohNLLc4WIypMM+3E/JWlX+WOYEVa7Kd0cGVrXZ3ROykLRo
Sld5t0W9VBGmQ9QCXNuhs4yjtN+5D1l0dEXZq2DhWC+5tQOOmOvzDytfzMziE4tpHtJDr5nCF4w4
hwXoDunz5rTKlpAhITyw9usESuH7MA8nj0RSZMB4LFXvknbBzjC6i9mfOqM7UpM/hQrF2SbKEgaF
MbvmAE7aL0DYmVjxhGzFwjmnEB96bMISXuAM9co0zwW83AZJX1MOZGACY2hOWim+a2bVom/KfZvG
3+JwmPirbL7xqE0sTXTI4Aez6/haRd4xwCxS/XQhZhShyJpUqGnHI9ZkhkiVwUyhC00YoS1sMELl
G9AZFnbLLZHBU1wrRvTNnniJZyAt82Sz47HpnkqIiF931wlLLjCKWbMUarc+8JrFgadHfxvosOMy
eM1heqKaqfUnEsO24S97DqTd6TXTCyZGTGpdE3RV8fyohRxGDWQaILHg97emaHz1AGDOfOSQUMtg
R4gcd32R1dCkHlNBDROw7gvL9nQ+mqlFpz/bn82n2X9p5S7s1c0xqGDAi9wibQAzkP0DSeV6/hHX
Ui4AERIHEvLNAbQOnhpuSo+0LygY3nXuKMIGN++cbEhMk09PqOP4/M01y53onl2lVwSpFaX6AcV9
l0N7VVFz1Vd7iGb3rNuz6fZG1JzXFBOQoFVsTI+rPX59hBH/RZrVDkan792hicg86U0xG0jF7vSL
gzy60WRbdcAThmOU6YCrwRZLZL5wk9dAQTc4TIsTl7n+Mu6iSnCDmaRbLrU3sW1zxI4r22WvGM7z
m9XeNXhRy36RYf76em+qqHMHqjpqIL4yvtmR5vn5d67smk/WzmE4TfmlVhF5zClQZzPJUJP/61ed
21TYV9apJVcqe2Im3ku7WJHfxzeXGNs0t7CfyqpG4YF8j5SjRmSZKs0CtNal10H1Edp3Y59jxHBN
TBqEItK4IEmrgeT7h+zK5tgmrvAz2tVxn4oh1a0GkXpdAyQipFvuiaN8SJcL2NQZa0BEn57K75Fr
S4gfuXd4uHNsAYW6d3z/VgVt+ZnDUzCFU9DnqFHTvpGxXZ0aNxAY0yOIg+Fd67P61n0OebqY/XC6
SHlyDAiBD6wX7Cn0k/+Fev7qcu5+QSLU58RVX/UP3oz1bUF5KN4VfUPR8QLesoy2CgkzIfXGygsc
RcxbkF5gWyC57jboJzUG93opvr7g4Nn1kix9xvBNqL+fWPs/uUJeMgY2R+yqY9r8SAY/1+/TpSEP
fwTI7t79fU4175AO7R2IvAzMO8emEK/yujTOC4zLmK6FJX1bq8/zGXacSJ/+C67Lj5+IYDdMCzzQ
sRLtdB5WskcyfnrFV8I5HolVc43/8RVv4wKTYHQMgDodAdEsjf9sOJtwpf1oYovTga5xoT6LyAPQ
3CILRqRL9ZMuFpsxxjVp1ekBJNWQXM3k4x+BPr1JsgJUV4QtUHRXcJC8Y5LMpvaZZOVnfC4yfAiO
EBl2Mq+Rle6LSBhffeaXGw+EVVt4gUDmjpFk5VyuKLRP/ZGl2eiW+hDV4GxLj9l95IOHjCqGI109
jm26jswFeXcFDTuEgF5ryHDrpHTcHWElyzrg48OZC7hxuojPPGZidqXIzfd3KhiYFxrI74lRXHVO
oEWVMVS7HUyKlx7nq/yF5nqYPTVw8bUarvYqHHe6iYfvxjI3+dAdvYK+X/lKTnCXNj22fKiTAx63
dJhxJ//P04TUWoqc73kNbfXqvW5X5wRhwaugfZqUZEscNzZuyGEqR9RB+OZ1Tu6SqKSNRPFHo7Ah
0AEhPfaorzWv21SVZbALBTF9CDpflw5lkYWuSegIQGHyuZCN61oI6oV1tkajscw793/tQI/7VSP6
FzZ77UMx8+hgX/hYgwGrcL0YdUryAZ/tIiIOTNrcPlcsatAkRYszsJ7NoRdOpn4e7MXYsuwaIihN
LW7U0sthYSsZWHwyh2b47skUwaA+nh4VZQ1QNCFyW/xIPAIk78HNXrRIdteN8+i0U8gShSJwdNv8
bZgh4WGAcruMeMWfT8DrRQH8qPWUI+MjHCJpLER1InbL0Yfoqr8ZQO/A0LEHIwsNJFM1y0e6C0Lw
A2FE2nR7rYgEPDh1oLmviGV+ux1pAV8U75x4TEDOVa37DLOT4CREHEXsBe6yQO/iGLZc8Ej1JZSB
+V7OcFDXxbTp9ch9X0ipfx3eJSRAw/dSANDHIVfBnFaOdMqz1YbkbkyPais+Xg4xOXEJvovShB8A
lNbwofT8cDnIjutmUJr5Xeh2dPfr5n/jKislWAjZ4P/IjoE+ihQJ6lBx6zFPQF4lOxoyDOxvBfKF
IwSvJijMSVczllYg3rvQHIBD1Ts82l2AbV6FX852aZtLL3HzxuWOB4quFRjYzove0d5fTGYLU1va
GeDgC7f/4ch/mOde3OEqo8nasX8TH1BDaWiACOokyHWgSnkCl1gK9Mtsumq8HEbqK7iNWtgEGL99
E8YiHuwuVYk9K+htp2Fh8/6cFwELqoGkRdPc4iG3P9rODcJtmgweK0arOjNHZ+UFrSOK9H7NfPfU
S3y/gM8id+WEXM/GFFFQdlVvPcb9b9StCafTcEHRxrMBMuQCdiaW+jYyEmgbr6OgM8ODgAwpzpnW
jsqC80wtZ+gJIzcNLVfKthxp3/+kqW3nO7gzPAkEqNHFBfrLBoKKaL60gjk5rZzGKGGp2JEb+f8Q
MzIq3lP9Q2J5CwDNPJjTTV2ZPSVDD3W5ef35jLAB4sAtcRpnuZSGpWP9GXbeqr32M1Lw/negmIlg
uzRx+bXdZKizCTdrCFCIfg71EWt3e5Ptpwh6AaLV4XDKYNfWOqBvF1shEdxBzsq7jwqLRloOrHux
A7hwkRQViGMaH/tZRSAbtTkYDWwnmF7qjprombqkhyb01lx+IWSXblh9fAOWhN+4k2E4JaRgzG0e
WoV+YvDHLbyY3XR8/Qcgzr7Dt/bCBVRynT1tWI/ZMbPfdWNcWqhgJ0tIYtyuYArqrqSIyDSpCdbD
VbCxR+O6+BPJaGhXSwzu5a8FzErpzUBpVGPughrOsLzB80jtgBOsd3JufehWHR/NJKdYyHZSwMKj
yK8fSmsL3WIQ3HC8sPT83K2HuKGmx/roPzTjbVo+0ZmYU1v9Z5cwG0NTUTuMluiDZH7TVAcqQE3J
2OfP9TqZBJg36MYxxAlvNwm8OyixognZfjDZ2qFRe3h4H0DRwXngdAqbZ1ME+TU08HZaeL+r76Xf
dYhj6rZG0TsN5/NP96jMKHPC7VNJg/5t6KpCqmzpVH4MJKF0AugMu3PxxiWqYOXbXfAbakApdOjn
CUauANf3LXbQeK9JFJWayhkuGMl1wFNskhel3P2kNXuPs9ubrOGhZunMZCN/RV9XBdB/ySVhclP2
M8yiO4uPcSoPTSVRGn1Cz+wdhcvvZvkVsA8K2/zkyg7LxAi1Wgm2HHuvsh+FO/Eezq4grClVBNQn
udbrE4eq9JV5jWvn0jRKTyUD6m6gWd+GroOaWpeebCNa1x0dv/XIsFx3fBjdKCKu+v+wfbwedvpk
5zjxHHTydQwqgFSVq8g7cixsKGEzrXWXdMm26YHpFBbhEmqyggOB9aYTeb8VJGKd+5f8C3M4NeKN
T8BPeq6FyMd/cy/mKeg5IhxEI5C/is+okz0gLKmR7B+d+KD/CgbwleP+teLucaNapJ2PBf2mp6ne
q9FVJl7xmUOKgPvQzmuO9IWvSUQ4vPKU2gaq9o6tjDwqge6a3zjOgu85yVyPk2OzEdQrheiGrPrt
9KV7ZVgTkLUzpREdSIaiNz+wOB39Vbn1OR8Kg9kOiVyC6uJ/15eYRLjL8oJGNg4vrA1JvwkV5wYW
a6xEWna6durR64wJmChDOUhoNfpQ9sykuvPM+U4FjiXUE0plE0fq2zdkeFSH+CLnIMpoAdtb69ir
uIUkM41lfgPdgYqH2lyDa52x0kWQE25oDm/OSyDyYEr27kE2exae0ODzVgvMec+nR/V2xVJCx74r
VGgZ/pR/e6hcRZyXl3tslA8cEpD5FrD+yWEjfyKwWqp574q5XsW2nH+1VHXrMpgGQW3vNwD/mbQJ
0iEOsHezrzRk7QIlUbnIUDVWWkdtTo1c5qTKzi2tahgf4tSnsbeNO7oF8eRzVOBnfr18WB7Y4DlE
nVncaHyTBLOY2V74j1SJOgoIfJWT/JYBx6X9hx7RturhwcVcPebLj/DHHW5DxrcuI7JbtALvXp4q
/gBI6cTRvlDDZxDAVUtta2YsL5bbI6NaWHO3IQwvmpEOKeFyT+l/PPPNZi1t5qvH4Z0wTjkJVdCy
yZ20f4OfrUvn+7Ad9OeOL9EGOJpsXatpvkLVusTPwIvnlPybxayA5ujUfaLw00alRUqaZz1OV7Ly
RnZIoSiB2V+uMhpK5f47izR2bNAAKWsBJ965vyYPjLwvNHisBFQoiR29UwSWpuv7SPZ/A/PWvSCG
+VF1e05IucaTgQi7rO1Klj8Qkq+KRn17o0zCIaPqQVlkfxvp5qv/db6bdo78/FMeRiS3y44nMCYP
n+vrYbDb2HY5lj1nSOaqvlQUD2PNdlNCEhDQ1wZbNOU5ojoOBk1G2azWQ2c1PzOcr4YorztvWpB9
IduLhDYBo8YI042L6+1W+kDkKYfTkZI/Ief6Ahptoj2+uSgBgp3uDEgUE7H/zoSmZCsSm5mLzZ9x
zxeyxia6j9ahdFhDPHRRdkfZJCiDc3QVnG8G0+J5eAGiStbcH6EHvw+Gq97WDksso+Afs2Oeatcf
Y4rHGYmdm7iavzeUxI0k3mBfl2T98EuvsnT7wsJvHxQBsqodEAbFR/FR3tj1SXc6bqwQwFxnQGqc
iACU6Ofe4g7PGzm180cvxQmyH0PbHXodMkmHJNvRzt0cscjQP0a6NvlO8HUe15lZ6J1af2fA5U11
vKvgkjpaMoshWas4MdpS61Kn0w/rHg8FGS5PpA3TZK7oYVsRAZjlXLibthZKjrFsAAVf+Zeep8DQ
Smc10ZO1JanPuQUUKJGolV+C8teh295m0Gwdw7tSS0cOcmYP7FNJNnJ9i7qeqsJUrtvY73wjKzU6
Wdr/6DYhQarwYUaulFaiLKq/z64HFB9R3YlCepDlwLbgRI5ORfSsXLeClMCJn3cpmJEVv6x9XE1O
lOheO3rF1VrBIJzZU4dlTZKdmb9ARTYekjq6YIH4RpFQXBbjSXERml6TDdBLoCAxZHDMKwq5Zf++
e47VWHHTAlm15VJ4/BDwq84gtLPU2B7Yxc2/OIGxWMoZUeQFKSHodBTPaEJ3WTbrFEVhcEqDZSBX
DlD3ccfm2DjcDeAnC4uRxHlAa9rgrGtbpO5zH9t1k+Jk9oP3j0PxBiKjXWnj1PqOqlGbgd0X5ZGt
2ujEJD1V7+dOgwosgMHLQwuAo2Y5KC6tS/TBE1y4d1bYBN7NY584YY/VLAB4geoOvhkd0AFJ6g3/
uNkDTydk7jJwEZjZmhC1b2587bmkKj7BZCdtSanzAz2/0ukEi/aWVBXxyRNvcSXLcIqJpyVBemoW
BE3VS4tAu25a9nsZOfqBcaWFNn5mFqBQjAFaNRqeDAJiz6ygJijJ9C5cH2VnpkEZGDHtiJxH7g6O
keUE4BKUpi2zoOWmJysY4t9WpIgtShADmI1gmb3FH+ZPsoaQBWoRaTNBWbTHK29Sc9qDLRbONdxc
pnbqGh6YtoiAT8GSEfSS/JL1qlfST/bIRtBklWIK+bqD8DicWHTi5OqY9IJUrQAZAikS2pMu6y8q
cQbnRjoWLzRVEZtqrYPyYUFWiX8bFA0NLj3oLco7YC3hdnRrhH9hOiXe5jb10XjOo0FvpTcZs0bF
TeU/h5U1FeJG5eHmnrkjKZOPNwNluRlQcAdrUSaRz+0Ng/BkcOc86SnhcfhdQNM2VsJTsqJfNcPt
Y/elu+cRcGELlweMxqjyDEcAEWRCHtvFNReGh4NoZCVJObLM8qRrjrORFpF2BICTZFTlqiuHDKdA
KshdqYtdRVUi7g21VClS8qAP8fM+LaNE95c8cAaMlVL1kM1fJu+H9mtpMhOSEogw04Woqt+9yvA5
wMnyVilWbCwPEYWbOgm4DBPIcOSCfYeFJXwSztyM+r7NhraSjKYm3wDOAbeUDPmeaKgDaXPtY6Ta
57oka8JIhgEjl3ScszWRM9Cv7mTX6p5rrsLdm0ANXs7zcdYtLBMqbkKV+oSDIQEsDPYTzQXIY8SV
t71cwvd6yU0IzDwoF52nIpKMzNkmT2plBParm+dfKN3I242wgywoSCaecasEX8tAaz8Pod+sHeae
ZQ/e97fEZWUmdrHK5k40qeDJchB+CEDeQ4OlhI6FjPuPvM6p/6OD8uaQeJqZ2tzVuZmG2QXgEpgx
Dd2abnLjaVyvG1uf9xvZbRJMMiq7U4bSNJF+CAraBW78VMdAdVrnqReuCjFTD8lgtnpgKVY5ZPkx
drGNdCH82l/YZ32VA9jWAgF5EojVlbE6fhjcM5RSXxiCIvYS6E07/p5lZcRFVWyfyVWvofxWsFux
v6fR0RCjZIQpd19WTwGhX1RGl1iOOZrGMvl2dPO/yOhIcnNjXSifaoklVqHUmYrvhoy+zm9OiRyh
oV0CHrM8NqfmGvDn0MLh4xIbpyJ2xxOHTnSvC/S0NVgcTB6cHGL5wnJMUxOuKMVrMV0oJRfGz4hB
NYKJF0k/j7tdzas753u0x4XkwW4KaehLC3xUoStZ8fV3U6ooGXCBY9z7VpcL4o1Tljt2NHQ1hJut
lV82XF5vt37tlxTszB9K895wcGNWOJ66bdziEkoRNuZc2JNwJ8lEpGy8tiVo0m9/NhQh2S4OXGaN
YVhtGlYQO8iOxU6fJIuJLgH1ngXyeIgV+SpOxji/Xi7rQ46n6arWSmKGF0rA5EpLfOJAlqgR/2w8
BwCUnmtHsIJxJ+Tc2mSx/PmYzNzp0oN0cYs8GVPWRwvy+nadnKUNVVQ5FU0adNo98XlJExYjKvbB
uR+3IAOOHnq9fQ0S2YwARxFJD0XGN+UPkUpDYfwWRMPM158ZiLXRjLXrX96Yi9gPphkz/rWNQ77Q
h/zihaTZPbTHfuzIpTljDd2ikFrHNX5RToI03CJDmxC9qFcAq1YDB9qqoyDV4HKgMGsGhV9MpmrI
6OVr2+eshzIodgkOh2vjOA6zvb9fZa/5dZgMffJvRc+a1BoNFpJopPQmGFF24z2a7l/6zadwWU+I
sX4up/1MFPn6aEqWegiAf+PNzRCP8ZVh6n2fIM7QvX2FcA8X2PJ6kyxSxk+JQg3vjTQEjaJ28lDn
z8bVDn9ZGnwNnfg/1i2lQ0Iti5L8phj4w4qxeevah0TNKiYSQMusdF9WoBKJv6jJOF6uyr0YfwYm
m4AbCvo5dtTaXH8JsIYBsI5za8q8rg9h3sv3N7YOO4n8UUOjslTpWOolLkaDJpAy4qXxfNkFh2mV
B9XIsBHLTQUgEeSObV9Io5ZgONDyYX55s7AAdchSnnNRWWl9eSTNkd/a5A8JQwKbS/dyNes7KWdR
TIPNFB+X3IqBI2RGc+kGP0aSr6B4enrJUE6blRX2r/umINCQxyuM/qr+8q/lWl/ekteCrfIboq5g
IEzEfP+dfQFUOK5OJ0d1DJHlWW/hILllFaB8CcB8WRt0XFf38hZfWpKarli+JuT+NLG2mIucSdm7
yu1u4HSVYCK2emK6nwAXxgvr3+umpXYVb5EbvQMpFeFrE097FDcT4YDkGj4raltOFwlMmioa4LMd
GRMNlFT7Fe77Qqz1L7Tzv15I0wbp/UiTQ6DuYnw2HsMlxAtjjI/nx+5PqsMzrH5i13IFs0h7qJcA
fdKFvctNXk0rHKFyguoXjWVS4kwo1cCaBhHZu5859tvKEQ6Kxi/yAWVX85dy0poFSc65UO93CrcW
D6jxyGQoL51QZbFiSknrdO4Y53o8aAkrWbR6zL1nk22e9tcqRlYHadragPpNZaaxGiTn1+RqbzWZ
pvQh+AMYnF2BRMxPczT9Sk+VJrJNT0iQcEw9DwjeHuwKMf98I8PF73CgOueSsMCmQJiQcGJtSaOr
lFCCKgEbzxCdYU2NTRyp+wVvI40GOKU/rxtA6AtWXORjb1rKDanTybelKRzwXfnlOvrOhPbJcE5d
hjNz1tRg1Az5GNyuerdbIDkdB5AbPunk3NzfG/WNll633F+W6putRCc4Wth2rEeLO/ukvkKWfrR6
nwuT5Lz7SKOj9fGmQi5oA2xq8fm+s62gq/bKVC6jr1276bMl2bQo8kCvJzU+VFHq84j+kWb5ZFiS
AJdZFuPuREWTEvolZEvJGBYMuQJ3cQ1a3M9MJoEcN8h6MVppk4v3ztoEDPb0P0YI13eakHL3BuU+
xYnlZjiwDPtUU41kV/Svb6onU+1Kb1cNkVSsHtWyP1VuTBmTVQDMy3CHEH88IbgPwsgiDuGRcM7D
fymvAIeaKqHZfUnYtr1G1YmU8jojN+NIQqT4w0ErQ7TbrPuM1vLo6S09cIMXGn6xm0DWb7lJGKZ7
h+gTBAG1SAyzO7PAR/bWsJ687EbMjCAJbfQWMzoiYor2KpnHcwCsYILo7u0kVW99d9slkKm784aN
/kZM2jh/7EtVGnqoiBrVtuIb1begDumD5sHTXx44oNyZnBhiG8ndKmescdeY8G+e6OMZpXvAS+sx
n5WLZC1crR6OspraT5Ya7t7g/fiEkoogSglZzHN1AwUBrTWg3EEMrMRnmLnw1xvStKYAovbVXB/3
9zF0fs5jNQpTH3FsWZF2K4klWBxyXm06Ya9NifdLWwgQl3eg6w76cZO7siBOEAFMVbf4j9cTQzd1
ouKhi902z0qT7KBNoJxFKsARs91wJWAUuEJFnV7Sw75UO6H02T3s5/yhXDg+TECEt7v/kFvWl+Gd
iqbPvBlfKOT/5UFtN0oKfgIBLWI02cmg3fHlrj5YoAdp2RDpAREi0n7lAWtqA9fOkmSZLZR5xed2
wEZLL6NC90qn1Z4y/KG9+tuSvH/NbtzPPW0s/ho440HQOXKfXpNzQBPXo3a6s/xDSack4zkMesuZ
jAWDRIu+Y7DzoDR26uViw9/wMfD9J9AsPBaJt5AjmC3OheheNCZWC8ch6zFv0b1JA4gzrLrGZ086
EiY4KOBi1CTst9w+1JDeVO4c3LSxEYZs26/DT9YlKqcs5g+LCpXAabci9g38Y+Cug/oRX3JBUjCF
Z44Pep0ar7r6wbB6KnQRhsqs5mEs0OFVpYy5PfNNokJXUevYEoLPpUersXGUIlg2XiAe256+rkvA
rz1dSOeh5sJeXgapjBfv7x5cZO06LFfC6fzJEiMuUiQ/SEGdB59XUWYIfeyf19cU+PTuRXuK92xa
kXAyqxsEDhQdYsgdd/7t3nyo3BxHE0nYCO6bumG2jZ4dEhbIqim2ejDJUmqh8GKb14IzpTQh4OJM
oHIIAQjyQkSn/d4GZZhroX0fvOrfIL91rCIJX5YfCiMQfYrDNSOJIIV0BFz2c30u0ZOPGt08OXJh
Sc0PAR/1Hm17foSyX63nW2GfZc4vUaPDzi/gJVIxJ7urCZJTIsQHhaHy1wrzSy4EYn9YtfmzUKIt
8DGj6akJ8WYFNH90fBawRiEnhbG6KkHysatdzc0pgNTiHXG69yfl1O+c9gMtTPGfVw7owsAk5Wjv
QBRaAfCF3ho7bAR9fDMBAqEmME8yFOYk69itEC4L4DvI8roCWKLfRMsex6a/CfW4QCDv/nJZKlZm
zu7CsRKe4koekXnxHU6Y++FtZZBaGvdkQlADORzS2ciZuvx3hf1tQZIZr+BYE0xsIqm5bBZFdPLK
p71xNZXXuletuYUO03XCDgHX15uwRg72euAqedJBupX226l95qjG6UxYNy2sIfp9Eq23qKAEsIHc
RuVJrSp/YmJ0ftkOcFdE48+qbVk4Y0SGQOt9VjUN5JOq/eIXhrxrXQeWgdYknHo2eBEeu6eM5Caf
sfD1l5bGBmTKFH35BBKr4bjApspj487EhR1ebQZHg+khr03W85zxs6wM0GfAO6QF3Ag9B6Ah4bDV
IMesgS/Porai/k3WVkKnETWpveb/F4gBDF5RcA0js/NGpCXoUs6p+AliiGu02XT4EkjiXBZnD5l8
Os6mZa4P77wmQBJSjYyz9Qy0AYM3sI3xCm2xXoOke4W3z5RLJ9D491G/DAYWG9rtecNiTxknEIP9
ef4GzZ2eJHC/N4BmqRNNhEH4xymCb2VwSdL4UrX7wMrKZQOggGaJRHoRwhQN80IZmjD4vTf7SNZA
OYQOQFaCSnS/75EIFSVLQiwsfszmmnf3yqBXtvylLlT+lI+jH+LwlfoX6EN04+26AoR5o0vcqUbG
PYeGmXCuj+r2/Nctns5E0TqAsJRhaMCccrr0laHIZXdtu8ZLswTaohG0JV80oRnuS3JSqq4jvxYe
EEW1RRAF9ShR/p42O2wpwWQruQNlNh9g/FAgVGJYrMlaVzUtC0xGZr1iyFMgCYXoOaOUZ450Hoj3
4grxH79e7yCgq1hPHIII843qpEKFt+5P8zbSpcJDPSevVqbpNHduI2bo9iAIkMuWYDdewDozpOio
bRFG3jVrrIXQk+ocscgVX7hLJQkoMylpGxwPdIby4iK0d3tlzEKjhOnXnPlQWr3ZVOhmhxzdvPqj
SDWCvQlvmgyE5k2kfKZS3EVX8dxAxgGnefu+3xn1DV19GobWKTALu9cdpigDd6jp5OiLh60/eoch
5VwNqVAzdESRhmT5wkM8xi/C+Y4s5FqQSXyaNVr0DsbH7u9/+hzTntwJ5qAJ4ultrJHak4e58Izy
v2IUpDW9sgTytXvYVqUXifGBUvn7oL+/akt1EtxHnSqhpCxIGFXPnUaFl0VAOYTGn5/Y4nFO4l4Y
XKeXwfVEDJfZWg9NiK8qyFZx5pCQ6nu2NELWf+XmZYtUiDbMIrvGb3FEIVIXHdlr8KqyB/XmTMuW
AES7qZ9hed3o+iMQk+oCTLzZuJg32qot9v5RbWeSZ2eSWDrcxNRTpKGuMYBlZaYDPT0k7k2c7cXW
1Dpy9vPuQon4buKkZts2tzeJA76jeZ3xe5noJXqPbp4dMHEjNQmpOtmrOEWC8WcZanfppxcAM+vR
Al727paTuX1NA9gfyvwbwW8J5H37/HyyeF2cyTG1mCzf/QtFWJiP0FIbdEB87Qh/xAFrR+mHXZH4
slrEAmeMYzOJHTbM4PW1pI306FiQ6mvs0udjPiWRpnRFji+wJ8fYiMINN8LzDG2aa1Q/4x+3mxPu
FfdbfRatl28FCi8tpogpIH0wPucxafyg+DX4zNpUtuzLWtmT3YvE1XsmKs4tYOfQ0o2Q6gEuCwhi
Z9lmD3JoQUpwNiFJYpZQkDJRPEQ08YuJ7g/Kj99sUfs1jQ8ViHojkPpCK8sJb/uWxbc7TrLetd3u
6QoVvlLQCzEEdDMDN5044GdAdvdzRsXYP5aUFpZM4tCk62Xg1JJjSA1BOMrjmQLy9+5AiPFagzJs
oaseXkMtLaj/23A9153V0zZgRkUPBglYFYGQm2upFcYG9BroafeLLbnF1I+SD89O9Yg6tcXl/JFd
N1iCLwa3VpET4RKuobuVEUw+/C4DYWqLhMJjOoNTlqxTtgRxjG/s0dSa1Ehn9tOEGBhAB24nqhKk
sXG+vL0yZdVQjLg5innMXwgDOfWT3G9hOg3pQtaQKNqiGP9x2DRLH/YI4Ufn3DfGgYLacyWJkkDy
EP0ej/9rFY02pvIjYxX9t8dBxzIWcYa5JGG1v8d2h9U78AhP3lKkff9PEsB14gJXaemq6NS4835i
T9wUGE9gvfyysTAOMktGbqvwZ0WCzNtsdptO6IN5dxY0fKLkaLAWqu8h7vtE8YZxGpbsQWDD7gAd
ufj56gstgV7nG1DRVeKQEq6/GN1kUC+rwZNCuOJ9N2UxK+mTt/LikSCcYsd1b1IoAH/d7POA76PA
PMDBAn1HXWdUNznpWNLXUX0UboqTm5RmT6g8ASexIMhg9yAF1NW99GcwQg8glfEA/yGYwisW+nT+
fMbl+zIUD3YC6amgHwhC/E01pLbCJq0Oa4IQYoO99ZR2fHeqOhgYhxzF49eCV/4qe9tSeJRx6cXm
oFkMcNu5EKPYEcstGSRcykmcnRMltmIcctAQbUr+hrW2okEWyfiRJaQc/D4yL3YcVHl5ppnNmoMS
RrnhvSgmx5r90vXDwzpRb5akxDtWcaft3asNscUfGC45vruT+7YLyDjb6W+k/Xq14lCbz5JR+SfE
dGrIp3pijrPekHoyIhuRER8Der0qrJZXyHxutp54tRnXZ0seCqBHUBz6Sh3ilFI5SmCEqyea1sC4
BvgEWkU9TIW8aUFQkUO5msGEm3ag34NHyo7BQqKfDFkDaIPmFYfgDhELpk2Nr3dQIkDo9ZI9ya8d
QtqeJ7KAmT9QjHxDxYybRtcsyPM3eplteX5e+T4F0EpuRPX2vexfI2NOa1JHZ3ahL2Ad440xhaV/
5Con/Dd8ZAQ0hS3s5fdyaA5WhLvOMJv0zZKOzYjyhFg44DDZQIocMvPWXd1sqy5KcOgMZTYAn00X
FUpeLWfBczk7s4KESmQEaamiPAII18i1RVUWQvRiHYcLFEshd2Fz78DMb5plvPoL3jk9hYtdhCVl
dSQTUeWI+8j6cUgK2S8piNFXgFx6Johs8nsCjokAgSAUC9V/oQEmIec25OBxsw/XFqYsqsgiDiSy
wpgI5KERPUJvaJywQLpdVPMQpfeiwQPO+khW6yJkQBy451j7fASM+m/b+KJP4LHpnn9d3lP+/lx+
PDXX1irDQpA33DAY4OFEvm8HK23gPA0heq1koIUJx/WTxmjgjp/iDDmZo472iN7QPtNj/6slYylA
GqAGp1M+SiRVhxcSmeFp7l9ZXG8GvXiJZJf/TpPmz9IMOJ3YEA0EAByHumQICtZ7TJ5zEKrm2vkI
pjf5eN9vx25T+1MaNIyqRGOVY8nYC/TAIrdHxThD8f5SfaXE9sBU64/hxzVR9HAl+mf3AjuM0x5c
fXPi/qYNiyWfc9/kBR/oVZ0ZR63mS/zByHtyFM3GFSJ2m48oxFhtN3gyZBYb2xZG7ifOJf3qE7yG
KvU0OG1fs4nr08UAfFq/Cv7XnCPMFWqpCUVH+nEM4EbYi4yYd/u3lxAbErUuPxsGkEOuWGmQ+o5H
Gy474BAP4KAd5wy8luEFkb2i8t3erPOoAc/8D38ebrM9+sVBcJpoXTZ4tAK7vHJkwe4odbbN/6eC
rcf7c/DAWi7PATyF9jqrvOoJ7MFSmfk74O8ln7OzRFilPtAcBvlm9+K+e5CyuaWMd1zoGYVB7+fV
Lo0iGQwhtwmA0I1aJwXdvnlujkO3QEzHU0Dtng+DwLPsR6NnVS6kOV0Tx0p74qQdrC8bl8RlFiXH
t8xWrQ1KZi92C7zjPFuXdlnqvXFXNDZjLDvyS+xd6yfuCG1utPhL9YJPZPNUMlOr7gLelxAEW2Ux
gGjUjyOHSs3xJlv6qf2uSp3x84SCkkWj6fD1oeGxY3ODnlmCBrBo2U2/MMkNJ7Bwd3yZMWvfHrCb
2yDBQxkD2Jr+4ApYWnUv8JOg00v/eyNbWt5C1QvjdyS1ce/X1pSTQkbwLU3Uj+hzamVHn4j5dgDh
d+zLmGDhIukpGkvys7SxPzfjPNiw6Hb02icuHA7XJjW1da3c8Fsr31yKxg9lBM8KmOBupZq7/gC8
P3nkH9O9+bIsHSbCNLUPwuh6EqN2Qvhx6wFK2TzNZS6S2lmoQtW7w1nslalzgp5IiKT4zGktoWmo
q2h9QrTRYnsGLcS58iiLl6uMga7ZaeLU8RHlI6G/pmawLoVycUhX4YcqKb4vdohgTViba+w+nmIW
/1JG8CugE4NFtwusBLlPCAGBxd+WdscoyWAy9E/R4oKExmVH6O2DbH+2ijepSZeN3C0TAwnFUbJF
prqRH8XBFS4iauOpJgk6gEtOqGrG0+pd7qcKJlH6qrjRyxq93LK1Bvjf6jLGO/jo3LZm6aJ2TTbg
9tpDSRoweIVK47YpAunsIfhFC4pdnNwk8ijwFXsPXRpOKoJk6CDtUPABFD4uJ2EGy3j4SsIBJpKk
TfDT+hi99E33Z7giZV5W1muJcdYyzNqten+VjK3/WdDnGsAwpgWGrENT9NBKhCCNP9ZO7X0mv0Nr
9F5alHREeX4Cd4/xxEH+BFRA8o/jtvI3j8jUzROUKHFlqc73iOyHybilp22mUOM0e9Aeypr/kzxV
dqukFmNwb2soY6GHVUSf2YS09B93GLF3EblGxHRGYVZg4cCzBVCw00rHmtdIHMWaAv+yzQ8ZjeV3
M5efVj1hObx2+E70n2hF+aWHUa0CPgYj8CYyl5SElx0UkyAe/cct14n6WLldFzHoEQdIEW/tPM/8
Dgq0xVCG7Z46SaWJfbUJuBuTbg8nYNpPcjwUkVJGywXalr1ZYHu/1UFCe/+o/fjQJnoG+UZIlbUe
kJ8hpwZy7h6jWKl25k4zpYazPJ3XW++gp3wnPDVOYVoEJgkojlD2ekRy/o/xr85zomct0BplQssx
dzNrZV0kyK08rS2J19yVglaaGfhVpraPM9pCdDrMwFtzqGm8hsK5KrPx6/eKcWcTZQYvNUb0Xl6Q
37viPVLv2Fue0VyUXNrNArT7sKQhhWShzUR1xs3EeEMN/OoTHN5wS/OFmwTQ4vegmsICWZIx/WBn
LvwVTqvDvIYuYF+DGvpeCKe925G5yBEYmNelXHyPAV80pXMHclHsxz+PjIgPx9q2CYDo1F0NtkIY
OEmihjji/ZjxNrjaSX3vwZshI+dOQxBgq/e8oRRheWVfKTI2dCGRNuskqVRQDVgMNvHKzW1nbYMw
uQpyE+KufCfwQjEsjuoCa5cX1BMHxYUu4kLuwLXPTGdw4COu/BcretqFC4e7RYEBcwDqtDfls3qE
Vf7C3LjLMrMJIC5MIe0FpoaNOj9uOdofbQJNhn47u8xrK5kTUEKHDh5LGRR5NYIZk6doI1qePZpX
BCo/u4NP81cb7VT1Yg91aRZQYvpapniM6SNnrbAQ6hYxCccviQMsQkjtHrPuL9RDLAEueMjh3P5h
JezZrfstIjeGuUgwfQAFtvUL4S6hwH6s03cn5+nMAaHU18VP2Lh4/r/FJVYqML26fKlWB5deOhw5
gPn7/n0zjwgWjjERSfT6IPncI92ivdQ0n+/CaP8HzNOjskP37nsPk7uORiv5u6VBoA8zTcg7bKRV
HZYTrUtH3zvPTxdpjQ0bCrRTFp8NgAwu2OJCZEzU0QDpfFH9GsUxIwvkldrc1HVezTwZtpQUveh/
yioIMgrr5q4p5KrC2BVSLcKTAXEI3PfE464eGVi28g9a86mI2ZgzART3jz5WQXzUBDiOb/YrpHNh
8qAPkDj82TPR61eqB93tpJUd/0E7OEghDhOOtJXX+OpIrHnPHvqih9oVWHSDui0ZHuGu+oB6LnW1
4FxtUulHvRnso6fNH5C3YGS3zcaxCMxrqGk2xsufllniD8362X8Hd/rvuXsq+jEJ6tDLNjlZg7or
9qYWY79k+YSMt1L3PGVhK/7W6w75My18x4QxVJXGuZDUbM07TGNQMgZmxaJIcYsTPWWFVPzjYV5P
4Dlvnr64PJQHTipvmTSVm+z0Hf1IOPvihjH0TdiCqZr+rRF2or/p3yTh4seoNd5dPq2iUiS9Wg+a
l8k1uNF2S73UQ0Ggqf6kr6WzJck1ZdOWCm9HpHbJvrU31hC/vAMAUhNmnjPxI4+QP/oTwE0TIVDo
EQ44cpi40j5iqDEku9fQV4Cd8eVcb2z1xA+32I7TppCBOfbGeSXcOdYVwpePx8e+v2+npo0F7LTJ
Kw8yci8T5swxOEi0Sh05PgHaUqZGe7GNKzk2xVJw39i5QyMm2Quu957ejcPIJznk739c4qYroZL2
wWSvkl6cwzGOr8gM+5UDp72Q6uAG0wpBPr0IRz2g6bri5kfXVkq82HlwgILPq68WxjMwMIkHnNcV
dAa08vBSwoqQCDTuRQoNJnz/1v0L6KyEF1stCaOg6Y7iArwfLBrbRNNwjgWLEpClfkY2YXa1ZAW5
um4TKltbmy9LUhuqo1zZJSdYVRjb/QoLy0qBo7jxc9bXzB5vhh8bo0JZL1XBDHD5lJNinCLun49N
A+39PNo0uL0CY+hZiG3mKDj0cHbZeCA4VipGY7mjE3hASDlPd/dNsYfU4l5VgCt04nRnrDDE9ENK
bk/TuLsmyUH6vYpwVD8mDW5Vox8Wz3/H64Kpc0u5r8K8x496n0jsfk4uZi4LwxZirs8rFB12HYqI
2xDiBZX3qa29VbKiGC4NCQZE4x1a45f/6w5n/kgfbP7IptK665T+seZvAcGG9pYwQbqJ0vWSaAY4
hQ4/8ozrPai3kochNLInP7qsaT4SihIRyqDLj7uXUr4xo5su68TbctNNiVyqT35Ukxj3m1G5VNsC
Hlo6WT7qPwCZRQDcJbwGRcX8yBfye+J8FYaZMap2wvwEtEu1Iizv1APGZSG/3YcLtJseFU33eH+x
gJl6GsVnNUNld9DLZ53JcR0Ku6AXOkRpWEktdBQImDgkv/40aQUNZ86bybJNJhMKvPWyTjPp+OE9
0ODTSYcLzaqRX5N6QMUH6LevIlwDS6/X3+WEHA7vpBSrOnsq2yrM5c82bk+11dVaflCOHFWYoSU4
zYyPkRG1ngKCTuqJvVyknM90r2fsXyHWWrfEn6T4lOou5SjDb1hVunlMtFhgzr7RGlKn+uvDv8d6
W8bAS4+1BHichENPi3uKVpgPhVQzjd1Td54TqJf69hqyef4zwe6Tr9X2fxb916nSf0dsinYqIsdr
PLRLzqaX28mzB7GBEyYNLzJGlilsHfsvtpfNQx6IBdtKjESGilH1sRSZxS/+s3RPrWnudseDmtvn
rTJtzcoJnyxlHXKvtF/7F8QU2VfUUKe9UN8SKySgGh+HSkrEA+ChrTrDzf8BQlKs/BEjaiGfPtm1
ntmWfwuQDyN9kp4T7E0cEPFovk+OBfQj5Rvo21RQ+Bb6u6GTolvqzlkOwFVGiHWyMeGqgNBK5lon
G9VXzF9cB1jGPKBuJtr6ha9nQw1/lGDTAkgvfdChEKSfui8vc+fuAXibRLVJFUCVwsVL2WLgCyk1
OwdHcgtRbJmD5PXHulFpqdZcTa09agHMtdooXm1e+4GSyztzq0dVzOGxOJ4Fb6P3gpf+DP0Ylj+R
c8wExeqEk1Jc5W0VTtsfpbGvmufBB3l7sNvNMLkm1vqXWrUU0F6qRbX3D/C/2OwNvArF5GRVYc3F
pwYsW8UIjZNJObbC4omWfaBYjN+PkC3IyapvTFxKd2A5nfWwOQamLdFrerbWelfaUbzlNwYmORky
h+iQs1RHyWO1ATPxC56okW6OdZFK3dV43VC1+zA7LaNUy2BZWpK3PYk3REEpNqfkR9iXun+DQl9d
WTD76jfNGtQpIcLkHJG72tglfT7LOEnbnQR+GpkaY+CXhheK07h+5yV6exaI9OJgmg1fyEsU9qKC
A547Hhq9jHTUwuiTJjPUmHxqe3O3YqF6J2GxCplWbetfl1irTpxmxBOu2ZinIzj2UqzG6ty4zfZv
as4rdOZja8/b+Z3e+IlJCHfzbYBzDjx9GM6WRs5xH8BNzzGMwSwJaJ8sKbx3cr8kMvIMCaZKqewv
rP2jUgEhQTJbJpYJ8AMyldABYOjx/tcx0ZZKaItjZlSxTwNBKp/MQN1MUfUl1mtAIi+L4TtoZlIQ
6c4SsoEfv3P4ngLgVjSPxkXvwjs2PCK1xhgV/y1xRALAVbYhz8VoU2N0JGdq8FErZUZJdtAx0MbP
ns9x3gAo069ywpCriLyp56LPUjPQjFf7Hg6gv2doAjQ4dq8e0xSTUCXf4ZSyxg6wuzhNcUr8fz4q
81JEFLNNVHgM27AAAzhMsaq3LQmML3yz4T8AOL/+fJ7dAbiruSzC0jfgKiH5L8hGqLAGwx2ROEVB
m42nKKL5fUV1qCuPFbcXLRele6YMUKKDdkBcjt8r9g8ku67jADn5fqq5SWy6i527V7F5le4GbcB7
ZrZQ98kSFp1JFHDOJ9L7sRj1m3ufAl7rYdD9sdIGr6JgGgdn0l/d9NWGVPJarY0LcGNG+2ZuMlo9
CUFxJ5xYL0aIzThba7JjFlOIiXNjE28LVq17dTV2WurO7bXErh6jCB4NzaFVkt7je/tHMWbHJQUs
ZySOhcMBHfq/QjD23M0Fx30FeP/dNWwE/IGm2cCl0nIu9kdilFkO1Y0L5FBwcar/MyCJHQ5I62WA
QgvEMKxFGrucSy4Meu8baNbo1lE3Fkh6mZrKKVMeQFdvrjHbOkZyYsHZUl1nrpV4CfGBb5VVScbv
DPBHn+iyYF47oXqRKZbYC8gnVNnRbgcJT+pLLRX7Ib1hk35XX9KmoANoArxvZs5OmnGKbi588Lw7
/zMfg7JDfS+MVWRT9qmAFmF1dN4ol4FZmIKWjIR8W01y7X7wIfEYVgFUQbkVlt2vgrNPPb8qCi4z
RK1aLMgnpA/sx4lMprYm4bbLtN1uesZnXDbjL2rKJ/3bnGR3kElUp8YQ+Pb26F05NGGaKHiEnb5u
xw6q2ZDq7PIosJvl7LDpfVfX0KBijP6OeiKWHgcONTPkRccS1JtYqdsDRZH2RvtpK3G5ZZsRDpfm
CeAxoR6MGGcuFy/TEiBJJXvWOhemjqiqVlet0/Jf/7PiuagdhKWGbc/IG4mi69JhdAQM1mJMJDvp
K3dV+C69gWNorrqDayHH1dQvKoJNYMnuyMz+Vj5ZeFL1Vl4XlBc10m9QSDZiKZ5yHy7FLkEa4zpZ
/4ndLsFv93Qv0Nq9r5Ws9BsahdApZtoK8g7Ug3qM+QAhVArEWHO/fqs6QIzLGjR6cDWVnH3Il+Zk
DWjjBP8wAYvbTqiXO3g4j50C5YrMMJlhdbLV3d19IhAWJoGXyiiOaQe7Cvk5uuLHaJJjU+/5OKtT
eCFp95Bv0CxH6KXS5kg7d0hyj/b8HF4GUt7MZF6684Slgdb0/kSXKH6zg4L4/tz5EL6KIBbRcfEq
+bZwB6qKZ54LzYLIaamJSvRj7pktzPM28fgyrZbA0wqJwG9ShCGrxFFK5YsWDZYsK1tb0KuwSHhy
CG10cRxQLthEr/J+2hIx9+VkVptWcKLDj9SoZoo1kJDPuYy+pmwl9+j5gxdCZZ0Etq9fxy47EOG+
9yLMTfS0ArS6NFgnW38QxKgeNM5U6wCeQfVgsQT/dHfk1iK60l4IgaOyuuX8Gn89/Dw3dyxjh9+r
yKZoQqkC2MeaT62gHOTIODrr85E48w0hUdmm8WzCGoQZh3z6IA+zatoBGx+RxDc2CxYDUaGKmPrn
4NqM8BFY8sTYUiWpbw9IkY4Ruj6k0X6fiiK7KovHfpkc3YhDrXiYUwWGKrNogpYCJz47Dt2g5qQ6
Q4NCyBHYFgkf+tnTpBqxICJnIur7VvN/8WuJtR8MUnVArQz4BjuyGefHWTKOxJOU+BZXS6nzIMtp
LdRyeEJqzz+NqmXmOdgZUVO9/yuChKB4/VDcsnsMxWvZUnOr+uSN8oL02BIZPjoiX/toyGSS805n
oH9oSVORozupsfXyvGTIyBDZs4xk5yEcz6oCMafcxQK5TTbxsRtYQ33ConyjuvHl7zMzfjzzqWCc
o+YVuVIrUJgYjTVLapY7PizT1+Eto96OgFjcmt4KICibhCNo+F9Z9HtMUbJy/QFfC73FzEFD4c08
6mMBW/cmzFmtRLxXSR1a03bW2ROAohbtcX2pbPSjG1ooi6yDkQZWVK6IZotNWJlzrJdC9drJizeH
o2De5kBfpvKwNK+QMUwz0H+I7Wj25MKvoKqf4kxVPradVT7cHijOSKkKzgQYlbMLBkzwcqHj1WXt
K2VnoK27TDR6zHdPfGPyZUWG6el0J46y6aLZqPBA5C1g8DOd2e6CIgHCV1IKtoFK8yg18rHttB40
jb8rSlLz01BWm5X0jJux/IGn2W/2GCTUHZVakXiWcGGhnTDY6mF2Qmdh00L/TcW1NWipfZL4SRjN
pazTkqYdsOyMGzcHIPemXXsyJf1fpDPA5fkYM8jZyhtHiASe8vr9kvrFBVVz9oBy+xl4FYvmlyRr
mrcEWoIutJa3HjFgf3kC+RIdgQFp02NvHsyLb0KGfQOBWt8CQCKkYzqa06STUBgMCsF1SN/5QK6N
N1y6jteac3CngBacYlOlvDPSmwPuJagJ4vfMZOl8NOf68MlwFQvDT97ojhQ/1d0noY25elZfRDSj
n8cqyG6eIH6QPcraN0iCjP3R6NCGfOXhUSZljPcpT1Q/qCdjugBCGO1xilmqdmnhtklEdck/bGZm
01IE+igFTyN5VEBMNTwd4XfMSuVtU14iV5IFaX7zqMARIpB7fdoPgHQrm58kfRa1CI6xM97KzZho
KaLYpGumtz7hLVWSWwClSp5T11thz0hXT6SZVToZDPI4k2V1wpkRweSL240g9DZjcWW4D2j5BjJ2
ECzLLfUC4JkPyQdGT6F1e4QNDRaGWp3J5zGyk+2W69BkTyr2g0chTgZ0EtoPv9r1EshaAXrSCeVZ
ShE1EtG9UsWhDvkrjWKq6cFp4Gs2XGmn1hfZWF+wN2y5lzNW2l482huJoQ5YkGMZqg4AFXOQtHAD
bTEuU/HAWarYH6pUzZPNLPe6yuzScEmsA7jdHdz3KYtDWLXzh3i2iEHbAmlRKyYvEtPv+xJXG7R+
LWqpNoAdm35n5ejC9+oysPy8LUHhdWeZXF0kQ19x9hEcnDugqdJsxzRrzbXWpGE3IbVAH83Wscrg
5gZj/nq4H8B9Kud57KxYdZ3HZ0QexSt6vvSAx8jBWMm3zEz6wDc8PDMQ5BDRdDJjYc2wd4uYcBja
kMAcUlA+jjC/Y+gj2QBG+U4SM+gdYCC8j6/FeWbKCtdNCQS+M1rMPrI3Lh7LNckJ9cKXyrlYC9ad
2EjzAw2OKKiiDlEYuIy1KBJ9o50j04FUXsmhj3rWLWcz38swiw9dD9zVewC/XHyfVfsm6AqmiioI
Qre/nlLkZyfXuq0ldu7ZbyZwcu/4nUVOnt/RGMKlsohBFaNNQvHVDKXu4EaOYPBZH4FHOmBghR+F
Lz2HeR4ppk4pLD8PY7+OxEwdUYzHCeHMg4qI6q6ItFfhy7pcdMTykhYIFn91VvFx1Vtxc6DnylFm
ElzCcXmB5i7lQKpaL3+sbzn+Mv2gHLGczDbAwzz9b4flMiWbLs4zoZoYRe/OXEFcr8bSefvfVr+s
h8FzMql3mPIoTvSpYwJg+WtEgnl72BV3V7MoUoc1ewpQh/eiUo8stbvzPDDEVb9gOr7bBTTbWrNB
+CDqFjknHU0KZywoLR71Fwr3qM5szabkQvPTyayWcAnz7xKseCYFnzGj+IkhSiQw2f5CvS9vVZpS
787yuOPLWYjw1cfQp+KZpHvCV7YaJGDHrLQlQJqchqsqqBeoXcvLAK59a5dDD+DbB7UksHMcoOUF
xH6PHG3Jw+e4fFFjmYfGpJsQpgqfbyYKWltdUhi66yHnshJFT8KUgyZN5kfG1sYzZ9WPtIQmcBou
G9zuZFvoAV6/ErD3o6X4q+bsAWDreziiRa79WpgRr1JkWf0LP/eFQA/rG9LJ5FhPsKZ+rmkohfbu
MmIUsE2srvR8CIzIG5IcpuCRGiZicHT9X9if4RReB3gmCmj72koLpmy1uQ9Fjx8GIYxz2bJCZn4I
8OvWuS97+LwTsu0bs0DZa+Sh1MmHvGdVSfMK02fLD2bGiWyM1eUTDmjR2R61HQn0lekvZiG92Y3B
V0+FRpILla7XGaK6NgRxCii4doNWJX3oG4dGiwmnVVw/xiX1iS2nBJWRFaIGdnUuSkYWAXYp3YDi
cmo/JCrID/AaJD9SllRNHlCa+2XZCL2NjwtoWJKRKJQ0w3/Q73+v1FWV0hBWz5Y8pXntwvIJpAJt
g5B27U7X3BihwLIFydSUC4MzKS/LmRggnQfOfxifV+WAWfV6g1laQOt6EQwJl55JAP+jTwoynIGl
nzrtI5cLoizmHs7hNNeeT5UL3Z6FOj72aPTht2vIJK3RC/2J9qakdVGNsjBK6BkXE5bPNAtLtEYt
jjJ7Qej3mMd/9PqH3c4wybolbZNFukMjzlJzp5uTFTJqyqHsoUibFvG8QZMEdcT1C5HTtC16X5vU
vbx+EK/XJnVu2UrWmAs+GHtQpESabklIPjB4E2GMBVm4s0BwAveCRBB0GCEP0Rx6yV966LLn8qFy
yZ368rO+2/gq81zJznJTCrHTElB0XcIZQOSXcRKlq55bGNkXC4C8w/UVZ75sbtRT2ftKgop3IED2
sNi209AMfCEzVQmZEzGyrTaZkWAzsr94VuoQm0rMzpP0UXUcqBn0yuZkumwgnrDXss4WvFbDZVuT
MVlVoLh36J4dpEWINBHNPkDFdNcTTMAkS3zxqT6uzIQl73D1POxftGLDrm9vwSjFbJoTzXHYpxZH
pr7y3ywv883annEJHL6fyjjn9D4x3SaA7x5RLkO8QXQXWUPEY5EYvPT8x/z+VeirHEAXKku/7UaI
7wMRdOVeosE/erc7xCi4NhAstEoGgucIWXbaRiKqagHfHyYQFgSqy7/EoD2pxZX5Lt7ArLpJ6JJP
uRbCrQ1loZURmUSp4/FX7bzdzfcKdlI/7cSvPJ7GmM1esB6gh/Q6peyeAS3ARRy1M7IijABL49nG
R+ONVrpgaA/TrqKuIkVRgxmltcpfxyCBymYCNdmQk7o93PlurASWo2hG4qwHfScL72oapYMS5nG8
0vELZfK0MMEh+VHjAqksGT9HpRCc3unT1FIXv608jC3alyhkVXmZvRwFTsiGQyEcV+AFfQ9FzyJX
KccRyPPZR8kIwEUA7jQLZxfUPmlL7uuU1mP6JfNv8yImKTGD4UPx7iqWvrI5GVb5kK8csXBOXQwh
11oZXP6U/Rfd+tKQSu8oXtv3EvBVD5TwL+a3ZFyVUV9f+1XX5uqLVMnU+sho7PlbJkTF/vJOZS34
/uxAHEfAKN52Zkmza357TNTHQYtf2i6SfmyTjzF8ZTIYlm5fp/9VEzhNWmlwVRVzckQ5igVGD1nv
6wZghXqGN0/3KDjHWVyZQQFYHxrG++8/mw3QbBPVs1lZ/wf65cUaeiz9y/VBnIGjexbjOncm5QMd
NPA/PtuV9rwSWZI9ML+fYSeJsnOosNhbhADjzhUGcAHI16ov+fQyCglzPPMSz//rYKTPjaGzJYOX
KFo6UjJmisnldJSrZAl3rTZtmeqKxx1EmCTXvVrhOrRgMAggkz1Cy4jnyGBEFrMhG7oyFT3kSO6O
SMUg8DHBZUxTbIkPahRTg0mQ+XBXHmoD6bDbkdcIec2Dw0Sbnqeeaq0LezTObCQ981Fjnh/csa2b
3+pA9vJ/aBae/ZGQhW1enJNZwZ9LQi+84qGQnazRXAAg6TUMEV0xuqJRh/ycqXTL1WtVZivY2wuv
xeY0uyWwiba7vvw7ldDgQQ9X8o7KtQf/nkosGDsj/cI7aif172QiGMrsWihdW8/S2Ro/RKYxSBI7
BjZBCcsSUg5xSrCI2zaWR8Z0YAp2zHRMLmHw0azEiWxJFDaxBDFOilv+0T7fmCORNfTIx/h42RdX
mKNT9IIMV3X95MkM7wOa/UJy77xdKO8591z/8LVtbK/+0uf70LMiS388ufXSjivEcuu3OOIJZ2Q8
9MXyOXEVDZ4vmLstgpdetvYz3OnKaUmI/TKJ0FAsn8VWo/8SYGpTJdsAOf5cd8WMRFRDLXnKp7PS
7p5nWBq0qVin/l3sGoDp8uWXS8L8gGfS1v78f653WZK1l1s9YKnMZ1fSdRx6MDU+GVZUkmyT7RR1
sOkpqPyrA56oswPv5At0eA8H6LzQMuXDVMxmN6mkOwEz4TvuhCV857dE4Rd+OpnqkinwQ4LkLmpQ
F6o+5uKVN85TxjmcU2OIaktNxIx3tgK7KO/4sKHAYBHGloXElDTR8YGUjhMdFWO9X5PaMO5KPlHO
Y+CXjGF4r86HRSjRdsy2p54EN3ZVKBo7mHCy+VNOG1/F2OzVXDDGdF1TPyxUpv990rywunozAXI3
m51tUtQJSAJUrnY1KiZqHutVZ3uG+V/wnQalWUt5UnEaqNFjPixUfDLKEXLuaWJ6y+wSbLzPBD94
GceZgeG+Lu4qRq5fG62wZ+psFTQBgTyOKzU7Lmjj1tVW0aBX5rbXToa00eUEKCSSmjNf5azayMzt
V+FZ8JYHX1W2AJYD+W0iCYgsIM17zaigQH9nNfZ3uJVGwAnMm9friKHf4wgMGlZ20tLOJCRPxhwc
uwDCzXfMHWqgovBATpihf4JOLUPXyPjR4iOjcUZqluQ2jWvf0DwbG77ouPCTrc6j2dA5Bvswe54R
EofR3CNRnHhdgcv2Ige4LxGKYpCqtQLGIM53xeao8paoWAVjoRqE/uMAsbVfNa5Vn28o+huO5KBT
aqFTvvMeTTOxQaXEF/RBoECUWSnsawsqUfVegqrXAJCBcB5p8O53kKtkhxWcyplttVvld+Htcz87
j1j9JdgZEQMnbpx4hxaJJOwKPXTPzcGq/MZfMrjWx76vWSq86LWHT/R5ue7v5HQPPlEpIM1y7oqy
j6d8R3i6yZ7oZjloI8JBnPliB1Ckvh0v5gUHoUuSPDBBxX+jAkjECaLbjltKAxy5xmQJmyrOAyOa
VyMR9CzpoScpJG/T4KSQ1bdb4fEbH8ruw81pTmcse+dkcEK3UAZ6RPg2Xtyu98zDtjlvkTGxYCYo
eDRKguG5oXjB5zxpNwqS5Pz5c1xv4lZCp8JXyq1kvred5PnMzAIuQsbqG3UXms5L+1mMB60Inr1Q
tGXXEq0Vyw7epLU63sc4rvOkVUkbftgLOtHVkd8exZtYFFq9piJj0IKXCCoe4uKmH2s5ST9LrA/G
o3l2PRgYxHZdf6HrLFgiWUDgWl1PH+CMMGWEb6x38W7amTqEyMEMbQtJd4tBK5Jz6Z3focmEvIEA
TmGMdvA+9pg8fJzMeEhcQxhObgWJvJvKTi75v0XOu4AMCYLDZOKAPVyPWhQY7dgVHYPQrFpGjRYK
KYCz5feGGiGFBeJFqhoCX612yBpYEm3cUJ7b57nS5RMUfVQHcLrSDDsg/bxrpAgpBvhlgTXGbQYn
CwLF/4ROLzOYk+DwxvjhL4oWq3Eyd1N8B/hq7opzMf88x+cauLSkxMiUvA4/yea/OflpIS0BQjEI
jQWjBOjQfrOikkx9w2AdgOBZKOky+NKXpj4c4AY02otK7tGVkCHEvxIMujE3xaiSdRhMiPkEQ4k5
nY+eSM/6a3rouAnx5jSTUpNflHsmnXZaOdcsYuk7vwj03G0W87GUDMZWMxlF0SlQkUk0JkAM/8dL
5S+7u7tGyFb0hgTOsc6IRnAWspGWVk4BB0PXYVVncfrxlA5LjWtGlgV2zXS9QubgpeCJrPyER3jU
C8QUP//S14ckfX6fd4neyP9Hgk0T+skrP1xXHx30UJVIE+dKdxt4W6A9YOIJQIfJH7xwj+TlvMxB
3kl51y6lLaISy99Bgj5mHZF/EbEvI6vCfOZdRCCdPow8eIzCQ+M2yoIp9xEhnM0T3HkAcf3b2zzo
N5tV1lFPnHo7i2FOdUIdZHGk0O4ViIOqg8/LGxl+GNDB7DirbCRlJZyqst5MJDJZdpr/UK9YxDY9
ADyq2TkMC4Zv1ZLkwcLTGBlNUgrcwYpHH8EMYSyRV8VExzcL/5B6XWD3ptf+3u+a2ICSpl6uCwhY
p3fn6TRWlITkWHBspMOelIX4COG5fVSBri2k9zrVH/wo+cglGC2UtTwj4NkxsmgHqxPhV9a9I94g
FfwMfYsbGVzIi4ZzLKdZNrpPgTat/bLhKPXHg7as8+RqJ2vdTetHHdGToPCb5AEGw02sqOG6jG92
DWZ4uHg7k7z0QdHFdmhbkGUX5AWb1pCR0G6ZeCMkef3/ndZixnTU1QD4EhBkYmNje0TLc5W14Dj2
Pl9eS56NRb1PwXhYQileplvDr2//0+yGMfpextcT39BNl1Srmj0RwGxZhd9BzQOxXlT7+F6w1uQM
YBZlSGKlZT3MebhuhgwRYpBZEIpjVoUsP4YTTYFF5RGcOBCw6FBTqN830s7qtB7DYLTeYT+uGJFN
3SWU4bXE7b67HRCWGsZrLONNwtsHRxOrThIJ9bx1fn3t3JFw+uodTpH+pMPTQGo9RRV9XF9M3SBv
4ayH4gr3VujHYkxvpobslkBz1ILebaCNyQ+l8Orq6eKMq8Yt7uirgj2TbliA9MbywIk1Q81aeMQS
GN5g0t+aHGRM8cUvwBNZ8Jqt9V78jPI9qQ23qntfq9O4YRs1WjQwot4IQPh7Odig3OERhGW725oW
KLTLoSLeEaUTXZFv988KIdFqLVgycyphTySHTq9mMaAlxK2gjeip6O+w94ccfo3WKdu4YImJouaj
ql9+0iulx5jS6LPcab3AReBgioxQ2WHuJVX+rWAJuSYqTy4AmAJtGxSrobQLZKMLd1H3N+iPIlkg
hK3lCfKCE2cV7BNtoMKZowxO9AHAmMOQ22Pmoyhssh18Ghji0WqEk+0+ZhtDqU6QqDjjF6U4V9bk
mPvwdQy0glzPayn706Csc+XphjzhfItbywiRm0ezdJrPrfZk/lgCMmhl8ActSxlPybZ8l0w/t5Do
XtJ2RuXDwRwjStqC3MtKfR4lpyZM62xLoOMh7rGfFKBFsZvv5eoGrOdK9vz+SitndJbXBehqBiPO
xzWI4Z5wV8pYtn6nw4nTImSjJ0fzG7QICr8RWVYf6oNJAHZxm2DaBBzBca1uwWUb81dXR9SQeXB9
Rex0xo3fadBtjAkcCTk+nAkFOkAwVYJ9Tj+11zaCGskyC6xGvYnGXrq87m7jG99kiV6Mz4AbFMeq
nBjfjg3o+xuUDEHzFvMzDJ0spsD+UgDaK2mA2me+7lk3csZikQPF8zpT5i5+0Q/w/5olMgo/EuG5
9bEw7SeX1W/7/wrgJn+km5AQi7fnEddzEgqr7PbgTwAJXCqDLNlubPRXX5Azo9caFdJIN2Eyaqv4
t1+zESStFp4+TgPZAZa0FRFJQG58UZ6+Vr2qvAx65CSiOxvkUKXtejOLIXAHIs/cS1HKHYNA9h3u
IhTb9vlchlV3vyYXnM4GLUHtQZgBTE3tWq7VHQlpATY9JgU3pR/reYcK83xIRl+ncpOMr1l4+93j
hPYWH/I2pm+LcoFi5GmEQT3lLJHTUM7pzhxitOa2/00yA98W71SlBB735wrrKdcrTnP6yP0h60xX
Wsf0yHRheqdSXWomV7j+F1VFeByl3x9PIkbo/r5pYB9/GARbU/WfbSDJmjos4YR6bsy77GY8x+/H
PTdB5clXExCqaQ18iYJ7au8CnlfkWac9RdPWGB1wAJofAwuHNakLiON2CrSVaXqOCl280X4RLERU
y3Ubi7BCURB9mRB0zKM/EDo5EMy/qEITWwBQ2tZ3TKSIjlr2/CtSFucRVGMiPJ2f0Op0fT5ak2lQ
fuTtYSJiPnzSEg+raQo9twrufDtV1VmoCu9vxrQTd8q0xErpT/5+uWHw8A0LJvSaI20BU9+9gOlg
kYFNJLfK5mjT4MMdmJ95yNpnNkNLvQoKoQufocCMyySZ6dtgIit/eNa292Og81IWE1zHo96iX1WF
6GfB6Yo1be5LpEt6f7jjUGL4iJwCJWFff3QNx3ltbrXAMZXdYLyaF9nXoEGVdrTrZ2Bj7c+xhvSq
lhe2RWE7rOis9ZfQ1s3mkqzKH80qIGm8ek/ixXJktloqb0hrGjd8uPUfvd/EMLbA72TCuttJOIiu
AO+jqBdKaSc/SM9fSLCvZZDcRFeShdz5pvfeO32vayefXpYE7/ivVNQpz0BzJ4Md37gvq7cnDjF4
MPgugzsoIKVvs5/oIfV6zCDHXRvCwSobh6cn1NaXzKKOqDOgILPvdJ+A0MWj3T8+hCSetm9PNXxE
gCfig1BBF+BumoU7RTa9QEJeEWBPGJCQWnlkj6aWibRnj6hTXIQjGOQEEOEsznHhddpafHnxqzpN
hR6hvyJcFj4KdFM127skhDvsi7kjI0nK4WWzP1S9NktHmMIsVmxnVj7F2a4kUjZwmrd3JaUYweqq
LPTkm8v3gcPA1QmGaPM99a0JGswW3BvFt3JnKRJckPqzORa2zA1OUkLq0wsKiHzlBHla7hJZJUQ8
yclZctsnAZzqLF/7yzDcFWvBfAIUPzX5JwUfN7AuYuCvRvBnu3DSMj4iMqxiqZnP/I20OfloxVWo
0gWv33WgXGMPV47SPyo2t7/laz4bgr/TdOA0iuMN2ylvHR6JBhw7DrgULhTrdMrAWf5w+dBZN4EP
igF60cHyljjkuu+bgS5Ll+3CdYM5wIvPKn7K49835JQRem+dSS1KdUm2iudiugTs8PGpZhDXzca+
6XN+I7QlrXsSs9B38xMXDtwjCOlTIvC01ivUMABTHg4Pdk+KbMQX/PfyzJ07cTWqtj2SM0QjEsl5
hxPJD3XgmobEu1bPaWxnhGkDv/lvwalDHxaRUqnKDFv/jvoLe3fw+QhUtQ8tbb45rBkpqj0EYEnn
KP9J8hX9O54gy0HlKnpf8Rc2QEhUgNk/2rMHmmcCA64AyirRUjnYN5s1x+58HehQfYxIOegAaVc3
LiOIBf1FJ6WHYetZyks/gjbzSrq70Ai26jJFLnxqXsvG6A9bPnummah6lCORLmF2DDeSpPcGyCR2
XvQH4gToRPlishSmVlZr1SlfA7tX7MTga3H3/DUqxfW3z+iB0VtCvUDApVbxjZfwYhD+BdnOSwMl
dlr47zZ9eqz7ISF24y+6ayySFMyHKb9K7GyqAZJ2qj9oyuc/ERjbKoSjMYOmu3b2HIzDImgl+JCY
EdKcORgufkaOWVYkmQAj66YpUSPGZFNtOJJKCLRyITZDYMWv95vTXU0psLzx0fhwllkbXWohXtrP
HIwSGqJ9d/yr3XA1D7/wWiRcXVSSw5JWCumaXyOHd8gWA0005Ul1gID2tLalTviccsVsuatkkFs9
rz1B6yqle0QphT6FTbauGtfXMXGlKBza0NTa4PT7rrfCd+5tkOgTNUMM6H5+t7+JKhFiScsXb9ss
t6VdbuGx08vYawJVyvM7qXzaD0w06LLZlWLiCTQNH1NfqLPyKszBQ/jVre9o56pVKvJ243V/jYpX
i6N0y+rl2FiVUuHhtxQz3bgOEp6/O5hhIBnwCR1Msyl3eCahPq84O2S8JfWP6PB+dlMJCQ+Ik7i6
T4G9YKNnWfu+BuZIIInG+g+U1scl7dIbl6+9Cbtnd2knAJ+EvnK8hLlH51icMg/rGJDOpQqMJxrS
INcUY5IJmZA+yumiFDWD4eMlOv740zO3btOzv3b/LksRAh87rK3FMcMjP344f1O/O0kjY5t0qgSG
/9U8NGd9PHvPfQCTRDcPvDQm5BqzFMza8ZS3xP7Evov/nN9LZnZJBDGVC3i2EYqjm6B5KGKE9PB0
6K9URbWg8pRMqtiJSa5f1/nL4ZFHdJGkbD7jZmy4pUuWKbpw3tbDzjND+gTXDIJjHCezLm9IfD/6
EByqP5SjVRzBpaj0MRYYNLpMEpG46bP6O2kZjrnYASvtTWuNIVhTBzQz+dVqUmBv+25y0VNYgg2D
YFubem8pZewgZNGeq4sZ3dUKrCDuoX+seMlDVqQMypndpgx4TgVcN9uN+OEHhivNARrgApDXTYEA
LCzIegphxv3waUjWU7QoZNOk0TEbWLPKBhgeXFWJAS8vXxGGemyt3IuG7fHERJ45j1ugpakgOawV
eG2AaDhTB8CuU7Whulfdibq91xv9jtuXEp/voB6ey+GWzEIDzz65UjNMPGj7+Nyd8i5Q3dCGlRzJ
NaQ7tCLRMHd2VmeIhEdDIec9q7tHp5fQuQj56a4tPLU/1mtA2fmbbpkcO3BttpQadGANe1RxawCH
/wSUsJNi+mZpPV7+aJagbNSROKBAnQJ5/ga3uYkr4qBUF5VzS3kMWOtmOWSeOP7ngpQaByeIIz/L
YpYXYJu6JXHMbO/dKmEQTpPm4iapxRbEsljTFvOOQMRhdWLTYlHQRfPKn6g/+iGdzyeNHbYReqgy
miXPtEBrY+zNnJoCzkGN48o4tPeoAoiPVo11iTr/1MVZznz+FIeEEsXDXbsgc0MoaSlt5xfi1b4x
/dHvcrN2WobCoZoP3n3uhoFFAjkc6DYTRYzvD1lhYLy0WEOJrk4W9TAUX3DkuA4lZkGUu3eJH+tl
gY4auKKF3wtciPMprdV6AixhYfvpRisbjpgtrP4K5LVUV4PaIqweBJbWF8kgFGCjZcQ9wvEB8fUn
sHBtS3T2m62rdTkZlGAxT0mjpHU89hekxUMTdeZpvDxY1V9lExdYL+QfP49xctSsw+y2wOAdwRub
4iAq7aPixagV2+tasv0VAtdKOu7F11ZZTkrAmLpF5pKkUtIguls8pWWUCTIkV4UJtdFJOs45hZ3r
xZaRi3xg57Y5du4sceMgk0jJq41r7av1DorXjHJ+NtRXf7p53joZBfjU4NHU36j4FLy+mBtJtjrc
67KJNauzRl26zKLn0me0nq7CDjRCGWIKh4oAqP3hmKHJOCcCgs4oPGlA8v25kMWiC/fOF4jx7USh
yiN7ar+YJwTw3yHmORmo2zN3h6GZxSgesb5Ky5iOI6Gu26+yRYGNLLFbE78zAZMq0Kf707o3a+/P
6KoqeRKu98Qet9ocPJEpO7ZDWNFm36qEW5wxzaTJmtRQrWn+vtGBJxKKjpPPwUm3MiPYfDhn0v02
zxdwHs26s6f2a1Cm0ZEh31t9YY/pHEc/WUEQclQfKkxg79KpC2ZbQjlqBp/Paj9MXKMG7qRAmYTd
80412genzFt29qb+umjUOY6J3HBzeN/CxqxtQnT9J0AGnLcDI/3YaM579g7FyBMp/bxbP7FnEsH8
iWH1oFfCtnAlLUy2lcG1+7BhReFj0Fglyx6XoEdJ/jsdcWvfj9DUc3U9Ew+DMRh6HS2xPsEqK6Fv
xFCedWl1j8yUjfibEzIsISM1+Q8GSM2trY0wTVva9BAmBIMSw3xa6dLQcc70SwvKyaRjV65/JL5v
/yn2gRwkNOT9tKBu2Rlg7afxXa16VEYWJOkyLNVcv49Qblv4MY+5ico5VlmelGbpbAduv8cUXUXj
elfVjn8XUMolFPPOu8HAEgXkqAI5vDxKsbs2+2AvZYWFM5J5w8ZGQQyvCzQCbwnwAnEb2TzZuvB5
Y23j/fy29P9Y9Vy+F1onTamIMHRIpGJBeW6TUOh+RPLli3bNjd0vZHz5vosXb1ZYXVu8z76EnqZO
axsM9HmWkK4zpg+vfuJmf6OEEIgZya4JBlMMtOkx4n1jG+rdmZsCmVNs2ppl4tWV7zvlzX4Mr73I
6TlpZDpY0dh/3xJPj1LNdzroG32qqgqO7ZvYNmQnDxKRpF5Nv4AOR6J7YKAbPEbg2V5S14L0z6Tx
rGT+Oi/sWaS7uDMUfF/cUDuazeLI4ur4Q5WfehjsVkiDS7vzb5w/cNe0WrbLlKBf7Lbq9G7/3woC
EvmbfYwWdpPu3WCrC1DP0Cmt5syf2Eq9RhLCI+pOoJNGgGva5EEEiRmld/wOXmc3L5TUXnWIuJUt
wfe4VyaS7UHc7x5fra17LlNp1P29dT7eVr+M2qQf0Ae5fH83fiQhhnQAHeMH76cQbXeK0De8Q8zS
Q3aCdDsPRuGo1KOfXaeO9trIF6PT8gipJ2bx+R0TTQM6+WdhZqcweNfwRkhZ4OsTkwVNsaYDw43P
vY9oLqqD23dK3OM7zQVdtUSEX9zndsqC/2rM07M7jCFhTMvBHktYYYB0vm9B1Isvc/XbBptyAZOs
E9F2KB2/j1So1mVtxJd2TpSMYIPUBmLBTEC70vLZlLZe03tNLfzoZeR1V7qozWftFSdTeL1m75L2
smcb1f0n1z0V6uwymcYlBbNtM4i1cHFW9EX6jLQ4xf+6SPkITphT9oBSNiQJmIli+Pfi+MNSt8gp
Nhp0EXdHIufyC61O++OC/f8NwZ9dGPUIidXbEeXswt+nFKnAjm4tiCOy1wYOGOE4CKUIx7+VY8lD
S/t9YhOkPTIalZcDyM0oCS4uGAf+RQjzQTsBHU/oEa8DeewxQHPv7yy55MDflLk81VNot1tx4Bjp
MrhZjt95TE53/4bccOCetsHcEAI4G/dYLvCcZctsaXRA/CGvEic0tnSMrxAkHpKZ2lXPrnG9o/Y2
1QrQFEnGLFTQRmKP5ijkDw8R4bQVwX30IAD+daG5sF7eepBjhI7js/CbbrmL496AONVZ5J7zAEvJ
yB2zhXmniVE6IFOf5J5OrB0DCEvG3L0WFR5uzROCenNT6nsJvxpzlxrKbz+JidQ+AMvHfNxqtmvV
xEoFEAMLTIR/xhhGKKmDNjiceEzzD3GtG/oyJlMCo2b1zgba8zHE1OLS+uC+7p+Sl73aOrgnQRMo
FFsVxTn+vWEtwPlN0mm00poroNyd3DOSfnHmw31buimRXRlb4xXCLKYB60W8igglERZbwcgiLuV5
t4Sugku92qEuN3jwyiHxVhkwqIfpbiu2y3UwHHDqO4SDgquLFIh3xErUg83kPnDj570SGKhoU6T4
dY51DOFjBIUF98y1jydwXwlvEvtrb7Kq2XxY9W6i18Pq7IKblgbj0pKer0WE7MPq0iyK2PwE3Gfx
1Yx1BENbEF3OY1SWDpOz7AVR4dujjIISPI6WbJnP00Wbtb77rKiJs6BwF/xtBtr4+kuSLhYrj3Bq
VsXqUhlfBLkD30lgOsTfBS+X3lObEJ/tVDS0T7RZVUFuZOjZKRhVkZer15xNkGJdePvDl745DJS+
5rzEo24P71PmZNoF/dcwVD4D41+M86OkpMhRxYcdZjeIwlZK8RBDUe4tFrZJscHcbISnWxoY9X8T
EwAQ+Lm0pOzr7KRT6CKCoRF0J+CWIhqEeLp3OLxA5KN/A/+D/EIBfEJ95j8MGSgaMr47qsZXMasD
/1r79P73kwuJyp3nt6+A1RTx0kigDtGrgTt69xBnVXQQdXfKLqprqbTIx5nvNVplbDzHF+UelF5f
v8gWQf3jEJonIwlLik1OR+R88q5rs2KFnl3JUCprJhTylNO2gZ2TdECdd/3huMZyHw6KvFfG4COF
6NzY2N20Lv/I8RPGHHACJo9iaLq5DPXXLa2DH51ErGuI4XyEK+TlUCV9dZ5nhlx+RDDUAl9ph3zy
9tnuofKi/lLOsbTjC8Gpe5anc4nGrhlpShp156F88z4jNm8pxub3YVrOWvzW1mnohY6nOf17xvQA
8ORtKig2dmkhGfHOACadbR47PVMECD3ylak3tQX5OEwGI2iVM2pmcLbvntT8tocNB61u8EBcVLP4
EVL2WZO20X9BGuxWYeVxnx3+4ExaGO9F/5n8t02BY/LtGMI+Hxpgtit3pFTlGmFQuV/LuRAxzIVR
Q9Ewk+sN3pIX/373Fa9E7IS887dlDAIWORu0RNR/F7R1VNDlc/JlReGEeVgfrrT47Dzk988GYxPD
jRO5rS61pnTC0KKMGY/Tw+UhF94b4FhtFbscALQ+dF2VE5HbuejvuUjICdu5Ub0Oth3Q6uEcv5cC
lV3QU79+6i0233o80TxmC/0lTP6gYRtQSTGh64MfXY8NDH2baMivhvrUWAs6GKXhqm91wIAsaVJi
Nof2EA7Ygw0GOxtXcH8luo9WTSy6Ll7t7eMtcWT5jzMN4vdanWA//jSCEAU7gcCMnwfSyiJhd6pX
+71Yw7eS+0DsaAxJj4GZmY+d5gAeLZFoXXiKbKUQleBEURY4IwVpBrmS0EIVVVq94BX38aPSRVNS
O+WBjYruWFDQ8JXw0mrQh6+VyG6XM/g2XfH3Z4uL5Ghoyx3gGjLLiTy1cjm+8RI5m/2SgyRL8mT+
NYoBzMMndceJZdHx9hRHWYL++1G7e4MkeKJF0PqjrOfpKv6Yi9hrkp0svMyI5QZets1wQsuBUzrx
MCYSUoNIY8QfKFRO7wj2xkF/3wwwTZVR+4h5Q1zpubeQMaAhob0j6eoLq/sIXS9X7cIvYeZ4XVIN
um6fUsFa7mCzoUdV8hpmoUjtpxiW3XZDHDbTA57/GYU96qQb2w3vCaIky3UBtWoDQI4z2+cmFSvJ
VAVcFqF5agmwLxfTCBaydlK/ClvumSROsigvZPbDZYlgpnj7PrcW9xePmzfy+aahd6Cv8ZcpoGTs
WQzx/1bFz5pEYYETISXFxYQivVrWsZjounvKiGzJP31j+TCdGzxKIUf5WPCcC6zlt8XqDMUmbnXG
LNsJ7kCofHIVkotsVgrdX9+um36WsBusNSgFwkPTV2sHcszSlAYsubz5yckhpWFeejCLSULhu4PS
S2+Oe4X3zPOuMJGp0VSIOnc/BVTHFIi4dumuHBpEw5Ol8vZQ/pd38GnzXtp1uoGrwAn4p+g/oc7Y
eops6ryvh1WcZWAdC23QxGs6XZOtT3vQbvEnGSkMDGBh5cRVyEazpHBIbU3UFjcKzRKzueI+OWuC
ENm4IioqvmYMWHidMUqcqVsV18ivr3HArSF8gk7uHvb54XgzsLtGyazD8TrW/DAI6PEuZBKhFar9
NsGk5v5JOF9zFY3wR9FrcBETKXVFwK78ftNpfiMcXJBKISgEZ9NYsB5SCHlMprNlzguJtQlB2h1K
yWPJa4RNw/d6YvIeFMeh3J/o4+wkNuzJvCfm3d8kV5/Xg/ico0qK3Lb2xtPE0E989kvgKhg24tiD
lqFHItq4hlhhbJcwpEcUKw0GrQdWwsHnAiwAGEfU8PB1DXnrj+aihSjBJ+biKUFhHZ7I0fBcAQKq
6Z2DQYbP4O+/tBbfIubBVAFPGKeCsfxfwzuDGzRcXao3JBwudWGo6xmLEwFRF2lx2dAOBXNPDb14
RZwWc2ABLGcK+8k+Dv6EEcGxEjzkHxyDWDBFmzHmcDT8bWel4rVASyKFEsnjFoo5CI6E7/yeULZc
a/CzYOTeB/ZuxVESthL4zoy65vWNuXu/+Tq/vnYsV8XCVeMLZsIXyYmmt+r16t9hzWAnz8gT9oFq
cL/uHpjJvhGJiIgq52ZCAQ1fBfJtDXb+yfvqu6ykM0eNWu/ku9vn00bYgsei6wLeDaMTD3o0/JW1
TiJMzxGMVM/SS4NwQBlngyXD/3lhmrV0aAh7foQR/w0D0W41aveqawxSIn3Uo5IihJIHrN6thFeW
+3ger2YqDGyonGg3R1AQybtsDwOxMhD2CBW1Ax5rccAK7Vn+P1RXTjySI8+AAe4CW44zOs79kpjI
uGZ1y3m3elaXDu20akVOB0B5GrvUzqEqbGjD/7owoi4Ohkyy3l9rdABUnUYgwU7yXqDG3Nq/7Z1O
5VD7Y3onjK0Kjr7ySXWg+x4DGMnVoZyQa/YS/GrITlvOY7q4GSUzIqHryQComANgIWlwHRr39LOU
hPjNP3V6VoznULQBG391eGTjDkCL0+1HVU9qV8rX1A2zqfOQGmtJq8IER7GqOEiSiOOrCsDI9/w4
JPBe6rLqWw4UAuwXA/z5M2IbWiJivKXvEhqIBrPuH+B0hwBNA3qbRGG6jZvbT9S4naExUcznxg3z
81ZVZHZBTxt6h8AhHAKXrNetN4xZw1B6vbzShvimc/WXMax9DyvjnHq85g6zXxYgSB6nnDs/e2PD
VIoSyd1FeHV9cYzo1xr7sxITpI7/GrVA270OaiLJ6BpoXr90aVsoW1CqqKXI87Bi3qbP9qDy0xl0
GjYVTqFwOu/kGeHIbyPBo05AEcQ18Vt5OuaFl6TuNAF8JOTjbs3wpJQru5Z/2J7HpaVWy6H9x/qS
ezsBQjtKMeSS7gpmhetDOt1RSYVO7jhWb404IY8Mq2psky8nmXxaO8H8Dm5aCfbTellRdn7vL4Zz
pPJHWEYcs9RK1awsP+tdurwleASpNv1hgHY31jEZpu9z+QriQMTf4by9x4rdqhBX9XfcyA/ekHaN
QkjajMplz/gb/C833lLn6DoJsladZadfE+L0DCwB6rDN/qj/Or3+AwmHETLJyhc0OdFpz7RC9nUW
/sQbCm/vSEd/z22LjnHvOfTqAGgt9mUIy2U8bUR3j+2SjqXZzCN2w252chfUg+5mus07R8ZyscSd
gHG7uYwIdga2LfTXVBT4SBdmTDjt8xENtvT1bqSKOhELY9sD4UOvnpT87nDhXPJvQRLWpP7qmbOH
U3Z4/ZDaz3NdDovQXsD5HfQRR8Ej7aEPVerjmKXf6m1AqNrR5ym15wybcdnTs4pH8qy2FXLcIZ/j
umQ2cr3wuSv9wzfLf07llUnLt4eYfun2HevU4UI0kr6xDEQYejfl09k1/TzljEFGs1CtdbXecsrJ
+/qDTE3c6ZV0R5NYSn60Z4l6ldu0dliBWmDEkXQmzmxLK3oDBbV5ydx36SJAjuwfXKbSb+oFJOz3
tZ074IYFoq6LiNkIvjRj1eEYO7JjgaEXV3qSX36zo1b/5+22qi4Ql0ompud/iAK1wR0WZBMNu0yb
Kisn+gSmzV3W+QsDNm+ONSZ/l0QPdyJuyaWyD7ojqGWKtFHLgo8jL/Hv/3J9Nwvc5Sf6z/NAEjGH
he8ZFlyAEUgR+cTjHpmklX6+lt2JHOlmoklFas6cTra9IktNGcJ+qpQs8lgkeNG0GtiX/ba3WZh6
XiMCYNQvd2fFcEeAE7T2D5F5yeO40JiMzoG06TxLeAQbMFYDppKBN63NmlgslIbRFhCRDaZMtXwR
6AelPwpOot7uEt9pyNWBEp9lQqVDlycd0cLd1hlzUAsQHZ5vE4/AqlIv3s7TMFGsgk9XEGtVkLl9
5WOTGgXOttvpbxdT1TZvsAs77hVFvN96FONEHosZVWYI6UDwn9yIaEteO+tWycwbh1bbNON4aHx2
iPVc38I/CT3LQdRlCI2gNhXvh8mYEm+S8unlraBZsz1uqqCieMrxhCESBJU5/h2bO0RRMCliZrcU
Admk2iaqkTro8a7k8zGaalWbWgyiVMRhnFx/Jjp/5VqrdWWiqN9aATNoI7knccUuWDZgs/s05KWn
uYNrekZd5DzgyPBeFeoPCVKSbnbPCjYrmFO2oMs640oK8gYTPlsuiDuewp5LbY6VSi59cSWcOxTb
1gxlrM7qy013ZDBUsbVhqhO0sB0ZzepJKNO2Fx35IhkCW3vRhwQerqXEFhCX07wAgc8Xam2cFZod
WolvaRpYysRI7whBzroV5CBTumF8Ae3dPBmUG+WIPknzr+lgdrqhYt1xqU4TtSS3lYPgV1LvhJBv
5CjCcC0ZUEqwWULGMNIOxE7bqLMQCc9Dx785WOeBXuGCbXPfRUkOrvybCgopq7Dyt9PQqkaocP3I
765EYRhJ0RNhWp1BGJoIvxk7hNWXfg6n67EWorta6A2tL4aqw0/gPilA0eT2A6v53arJZ2ECzpE7
NefVk/YuyPq7JBSSM93KC9ni13rXZDgPSJTuyFqcmellMfavRduAKVDAPTt/GPPBhtE4MNrBs8+f
OG3t2cFql5LfY1IMCdWNmakwOZWD/Oj1jWNo/yBHpXy296mB76Hlq1/TzrFQEuWD/0/Pl2h+m/uf
4U4NgIWbYzmx4J9r9E6ePiu8O0bZGKSCmuVWKQ/yGFUr7Q/iBxR6cN3PuF1yIPyNj/+yWzeyZ6pP
9A1xAJetASGvA/r65sSehx3C+rzJbKZLpw2Y38Wvksjbxg19Wy2HuQzY5G4v+vRomP4MTzmXu1YB
YP9GB8Tmo/dgtuz1ed64P0HsWgsUdNgWESnC+ykyfwOP35rb9EQFj4VX9VFs3TikNXe4qPlDmLNA
iWSKRElY4BBUjiqo9z4Ag8ToX3LX0sMcgkXV11Vu2RFqM+b/oSE/8ReqV8tJAVS55JETvzVmFo0e
XLIP4VBXy6/Y9xil8NcS+plLSKysq3+A3U+dBC1A2hE1w1O6gcqI91Wo9aUUtQhpyRDpVo7+7i3V
xe8vYU/Fg4+Q+MzyT5GL4c+1hATyn7J/CMdzoaXBOzlMA5x/jtiexjqhvezAmuNUwVcjBkN3XkkO
y4eT6relhgHGyoT1ocFBhY2b03vteGOcgJzKa9Cz9uL8KC6bi7s/xcJMpAvJP3ubICR6ph+KPgKF
9HFac5mMW034tXI1mSc4xMi44wLY8Egb0t90ptYCxRCVOXnpev4NEd8L77nrmxPJdzbXHViUMHId
ulSvds3NCup42mJ2uSfvcp1Fy5cppsT6a2earUbO8DVN99rPd7vDGL0+zqzrCYPNlZ5gyLGo46rZ
SyilAiM6MeBWlxIw8aFA0Xbpj/misn2DyXmZBq/LF6hxSGVGsgiOzF8lEXxPf2aWUJ8XZjZd3+i5
6DyClz5as5lcFSnnqXmlVybI+kLBUejyIJ2UIFquvcLMRGAN07ihJTM21C6UP7rZ//CMZKsS0fvt
b8aq4GTz4vQXAA/fqNCFdQEl80K4/fvQGfYbpREmZRbZE9lcw6R64XO+Cl9MNFdqQGNHB5pqWazy
GODdQGteOaqVbUBSw2jl+yNseiFAghwNkP4K4TwMuHg3t162Nqswy/C3wMFAsf+lYc3P/gyzu6Ek
7X1QtSYTuEfxiDqsjosO1nohk+CSUX+Xn0+1IPqBL3IY9wmTA+XDoMSQm0fChaaM+0okTY09f4Xx
TNjUakf5aon+ooi1PfCjweLPWL9hAAtSwB/DILiKbGEuGgJe+g2fdQAJw/8OnFfOUs+IMiBG+YIG
h44W/NoQgdT+P257zOT/qyylVQZ6IB0MYHRFN93YbZiNCr2Ei/7khF1jeyYKd7LlNFTk05qWmHJD
0SyIkc9UQmOZFAoiMmULBr6CCBUBilI+xvEE956rAFH6y2zqy0/4/o9Ay9aran9bz7+QQwvFJ/By
pqvgCe8ewr5BNwmabaXnoDPTK3IuUw7XRSI2XbfTy+8CY8pcvmoiBgomulqkGuxSFczrmqc/mGm6
tviZ2PuX/VU9MGqPfLmRoZ091hELtI3pzJiSUk3WW+bpeE2lM5woNMQkum/2GqHi1cFIFqIAbecJ
LQSAlOmZ2yvI46G8nsJFPsZpqvoFVUUdMV9gjUp7ASaCgYb1KuvvESkcjFGgkuK7S2UhJY3hBnUp
qSanfd7AruGylr63lXe1wq7QtG7+3NxHMv5CQE9HfsJWEfsQfjHN4eq8+jWLdJcPm1/2JWDXesSY
pp2rf8RwxNyK7s9JLTGtKo+BuUK3SaQ0MuvZ6LvGufLE7M96P0jhBcR4OjHMN2hYsXNKOCRWtduX
uq81IapOZ224MvrE2zP2FEMWtTTSGIhN8RYJGppaKGZ0rERCkyeLh0gGaRqT9QaPhEN4AfiUe/XI
IIfDbfuG38YYiZBFrS9diitayCwS0l+VW5sKDFWBThAthBugrsKJzh/kQkIJKUJ2BKIi79/P9Uj0
Ir6pth7cZ0zRcrNdKGfQPtFHCKYTPZ5RJLw+xtuYEGRRxFYSMpeBlOFGFx5DheyHzsjktXn1+ElB
EmW1uVpFx4sSc1pBdkEjgnl83FtaMiGGGehMTiR+wuoFHGvLqt2z7NBFkiL65CY+KYAXMCmsXOVU
hYmGcwWxqYwmFB2tpnrFmjFtxztWqytSGJJE99cAtZwWUwF8jG3gn+j3HYnVXSI6Lf1wgc/yewOS
KXVRjmSjz1eZ+MEUUzA5zoKyACwqz39thYgcp83J9PtY+1dsoZ8uDkWoinIXU7ETbTH/Zwv0djEt
y5vV2ZOhKnoYIVZx62vNYOFzeVUsjQ5RBumMhnEeAYy4DjZPuGZW3wgn9ZIREFDD2TjYJa9/t0Sx
jxgXqD/lPx5cXjC+NADcDh0WdPd+8gR3UA0Hla1b/sNKnu4cHgOypbYwIIeyQdHk0PC+DYjVd/fT
A/o+t4XFC/po+wTJ+t2yX+q66Wz9l9XxFk+fbQD3N6p0PrLYB9i8BF/2+nZ9TvLmi5Y6VoCNZVc1
oqQI9t+UbqV/IOzOxMIFa1/Fy/M8SLPFWUhauy5FsxnYxqpL+KQdAGnihAbrGwDqo13FBmby37st
ANh/71AJm/Ig8UoKFvK8cOV50gkbVgFvKAS0asPmYscg4NgEqsa4VNnw8IY4cEA1/TDXyeBC8vxU
Z7UU5NxrJd0p40+03OgQJe95RtQL2odMb/+X0TPRRbZmnfi4NFz7BfCzuJ1O5x7eT2CIQax8+8Az
829Cx7+ezbxaxPJBU7WNMiO4A9SFf0W0zEbEChVTC4AO8Yd/qvwTN5WwY5xeWULdsWhZDbzaZMzo
+KCiGmTGfFvhtiX3ug4S0FzlOZwkcQ/7bdmrTBoA+sVeq3YVh+Rt2oZWO98KsOw7hOvGJqWsLh10
HLFd8/vczokaPlrO2AHENTOc0a5DSGzPbrpD7gFajHQxiA58E3IYARcuRjoySzXydvtSMYqJU/xA
P+e2tQCKnSSS2osyk2YCu9oxHoan7SDA8g9+hk0xzQpZ2ZbofKPRNFq9IqB0ISGAPApLCE90D34w
wXXo9JckAPIoDwd8MUhap9MWmE1nXgp9hLA3UR6kMu1tTdmBH7mjwf7hGU8Wzf8CKBUlhgXTS/0g
sumhIv5jj/89ldyRCiEwzjrx7vlISEy88XdnWRxvLSRiMIhKIY+65k+EcKb2kFyO3qaOYkA+LA5A
ZUFWH1Xmd59Zk/lVDZg7aNi9/7QxDyTQqGp6OQa6S93KybpXGpKVavkzMzye/OUM6HxDeQBR35Ac
lIwqpBq75qfFXz4N/NbgQCnW1hrd9Mqtq7xRepim/pPLhk8v7GwYHm1oQ0mzzuhbAuD0P+sS63M8
/EajaKEpDqdhB5s1IZ/477xFtYT93S3Z2ZrYIwzrSxEgrJeXjh5M4/o+UI/a8Va9HFy9Nua6rVWI
vupv20tb4Dms/IgraG4BLJhMtThFrD231+gkAcEvdXZ3DrQYPmkrSvm+c0wMCDStK9Ij1Xl2LXin
FjIRMsmS3nU1Tv2t/0CBYtTbz6/gH7v/EGBeiKDQRbVxuMjR3pThp8F5vHskbs87I83FAzkcItH8
MT5CbfBzTq7R/hfQ8m9VwFvy3tMpCXM8bTbKzs0A80iOeu477/jC04lcsyZaLWcbg6CW9mlcjKZ8
pwX+b5l7p54WJVWaWapgy769kXi/QfM+MY9oSF2F+z/Bm99ja4X5uKANw/qp7QxgTb/xdbYcg2IY
YFM9HnCTHUkk5sXmCipN5zc0EG6EUXSC6D5dB7x0SYwBhEMH+qLYyPXUe3pmb+NO5Qv+147bZTw2
3W/bI5Som3v7K3qSTE8Yxdkxbg/rUzStqkyzwJ3+HL+U1EeXdSKOW+4j49yZuOByhDXyZ54WnoK5
1mtGRP1CJ3HilxfQk6CTVT8NVxo6vuhFXdpIGqOn9hVsRcywM4rbHygcITEuQuI5EhEWFWLvfMGr
Sbd+wis1vbpAYQGXkbZlvLH5+a+HQnqZQUzTMOKv9wY/5HfHN6qlc3sNScfsGUhJopAIlHV/jggh
qNgUTKMm5F5QoYL0nGekgMT2XR7aQjBFc4/OHH2UQG2JZQlNm5lgVMWQWP9kwrLr0UkfP1rUq1kR
OX0kA4/7ELFBGFcnzBEUk2DG0AS0Y9bRxVyPHcGSJ710fE5fy0YsL6sMVkDcEYY5LoUjF4aVQi0G
ysAT2/c3w2mXiiLhUAvFUyEAX9MZhd6BZd8FH9RyKww0t6krIF36b7On2ZJR1v1GjQekRWDyxQ9z
YcgZwgROjReW+8OW4fZF69Xpc6CWpMUi5JWW3fyEPAERCo2tTDXxdQyDXa1QeHk1hM8gOXrRuHDS
HtkmJ41pxGZxRSroMmuthzY998bEbLoBLfO5XVa+LKc29xoZCf41JJ2GiRb4WSSaLYStlaXOzGfK
xkLgs6cn0GDaoXBPUYJXwYeTbGZGnmVqvDvFVy66l1VS/B/zyCEgO4zLZBE8G9mhNsiHNCmJT6dF
eB1FjrkbuxMLwnPwSpOEalaqRpeUUtWyyttH3blb2qF4i1TQvUzmR0ZMhULOWj9fr75YsLdZf5NZ
sCr7D3MDyAuBBkjRH4dfP5OuB55x+AXf5QaMNy6JeZuetcdiabQ7w0neayCf8vhqX8TAiOHpClXt
dku/eFJx6NiLp+4I+KLt+s988ymAy5CCgFQBHid287VcJRHS2GKtixgPUdbWn+8b/0+gYRik9zQI
QcJllmIadvtaoJf86RvMxle/8wOuc26+Ax1QLPpIgIlfZguWsUsMDEe3jA0dEA3NcfsHr2GGb6fy
Dg/i6S8njz/IvVPHIOZ4WqgeZmVuQWprZlUfZAblQpejR3tk62MCHO9hoLGvXyktF4FUa55J/cIg
Z4hwRhpH2qWZTEqeu15qeGJrBJaAAofx5EY07S79SKzU1ZDTvzBeoTpXuP7Cz8O9X50H6h1XLdyI
fdUAn9PqoNtK7zMD6plQfLrjhVyJ4tV6s//nGWTG6qt5/PN6dsekSJ1oRMbuDHGMpwZyZiJiVA+r
+Sz7IAf7reT1nhqv7qoGKFyjm/axz2SW/JvWXUhgxHcOglCsVlYmYfpDLOokKZnkhQ+vIVb5WIf3
M50V70uuYyGk3xBjgOSqWs7mQYLy0Z7XO9iBcOllRJtzeOSdhRFhAuyZ3+JQEKK4JihiwJenZn+N
5wVk2HqCB0Uy959zo+1iR1OXB0nRyouCNNSioONoB3RclZ2rBBWS4QRwab2keJ9BV/7c6o1qmxyG
quuWgqzFYpY+5H0DfA0Otx3AVRmeWYv/rSR3tnN/OGvXJbH6yPE/+bCaTusgYR8H9eC+hh4IIhB2
2Rzvv0dhTKqqi7ME/dxfTeOnhOeUws3CAsnMUN1wKWNNV0dwXg9Ip06WzToizbO3v41IRdCvfV8q
UsbFag4Bz5VjNAbbX3uuyH6bAappqWc6fiPalotkiVkAf4ULkEC0WGTg/3+Phclf+1+5G4Q2nW9C
01Sk3GL4AA1JNwWPf0Mhu0VioU86I4laJEmb58OpySabTCOcAGHOy4mLjyZRcTZj9o65iJXdLZ0b
IOET48Xmmd7uvcb5/7rF8lKUicsFl7SpLmzYJtbLH4jbVvTPEIupVo44VtPtlHMA6ypw7sVphlB1
0oMkuet+RVXjkceL4xI10C/ReQ+fWTwPWXQvsEd3+ra7P7HdTp3Qnfb+9NxcDH1JC7EQwPgv7baQ
JoXaNEf14ZawFIqCXlMaADkF41PBVmUMeTUzAGSxppCSu8PFoCgNok51oEUoQJVyQ1contpll6Xy
aGWF+SdEV5Tzu2rpGku1JndoOoN1k4kOBsSLRblCLpa+00SR2hhmirCUxgoYfEPMwU+qBQTsbwlw
HVMU/+GVYNKiHxCjhDRQm9pgPA0pkg4aCJkJxMynjJPCBNySyiD3rmzPtwnowvVaJSszPq569/sS
CAgTyvXUVoqgQpwITH7/oi7MyfMcLvolkPulPTLltfZQ9HY3cz+FcOD4/zzUBh5P8q+hwnSKnVeo
x3MPKvWvBGMYLqLuWsHdUU//TutsEfvD4KM7LfP/moygHItk8TzkPE5do+rcxxdKfv/ZFNre3jbU
arHPq6Sjv3JFyjVFT2NbqR6nmQ0UQ8VMCdAS2/jOSmUvgV0HNHczSbmmAwLiFgpowc3mKJ62YCNo
it0ndTCDlXSVxh2ZYwAjFWGteR28yiCLc9FAOFmmI4aQT5dLS7H4XVHqtWNXur+Dq/3ubCvFt7Ft
sKdxaA9LVUgEK0RhynkI6wx60gQkpTOYQFN1M3z0B+sUwc8q3AodF7FI7QUbrqFb9lPrtiAykF3p
nhZiervoq0ThbzfzmmHneZS8OlB/oguD4kPUnaIBGQxWeNVbGaGh7Gw3RfOfMcOMcwbEhmaEXHWY
cd+HBI7rwBR5lzwT+wlHT8Nsmc7HvwbwEnEbuiYcC3f1Ahe4y0j11lYWhOFmLbfyzOO12pUHheP6
vG783sDcZVMZZF5vgU2c8SiqXuNJ7UBsnd6qLNktMAzIp16wXtGYsYe8tSmBchKRtuH4mWNx4Q5c
m9gP+ZCDo4VuD80cjRpsKqGzVeO754iBo/03VaSruJ8AD/tD13cCCK89XDqPM/wsblVJeDu/wLxP
Zl2gMB/bAAasxs6ZTpXWCZxQ9cmv9bSXb7jeWT8RrYN8saULc/MyEeglgEI00VcpNYwzzJkMMKNI
c/QKel76+wut9JkJy8hqHXCTQ3imxKx+7lYnIBnX8OZrnbt6TQGGWM6X9kQKNqdtIsK8GthsAjgA
/kaMqjw0lCbeSNTW5MLNT0e5RmVSp54v/CKFw3irA6ih0xotsAUmUSVUWaetvgKY8zEeplAp6FcT
K50TnM/ekjbn/ywbJ+zV6qCRXWC7/fWoy3Ojbl+HExvDk/bfNM90A1ZyOIY5jkJnQVl1GSwhdmaD
2tXp727Y3PNKCc68OFei1Ru7lAdJxw0fhZbaBM6SlG8rGZPCccFpHiyP73sllEYTtTaPne7sgD88
Am2DbeepMXifG65ruFxLKeDEgIxzP/bfjuzXBhEN3ZDw/n1Q0xtFOR3Q9BvMCtoaOgpHbSDqupoW
rIaLcwRo/RBraorBvyiJB655spVHs4LYfLfgymF7zcXOLW9YHyuwyE6rx3ENvMwDYRw9RcdwkQxi
22SytY1Kj2fZ0ofZHbKT5UTZQdVjWYdGUBJg/uLdwSycU00tn0Ioc0VfbcLGylv2e16d4Lf0bK+p
9O+kahh0PR18SW9DCM1TXJzcJxT+fNNK1F5BtjQ9iv6samuRRqvgzNdCNBJNALNhThqHH3K5l9wS
+qKjhMO0MrZXQh82spOqUek7apyM+kLo10nqT07plpDefjzpgWGQqFAcbeYyRSiSlj2BhqBCwsf2
zuEI3pD6GRIM7Kg7njhF8VbIaUx+mkmO1iBQ+cDMdXHwENK8+JDtB4kjZSWPTgGcbmeRApZITyma
kZP1p154VtUquVSdABuh/YdQJBCA+Ev4BK+Exxn/2CD2dMDUwriHE4/O/Nq3nlCvnQvMZ/OxkQFQ
hOnQ1fzKD1BMDa6noU0Qtevbs4GGNCG7Hm/F/1cAED/CrV2kEhsYOehRH/N3HaL1sGaDPHFo8YLX
IH6VhSiVx5EkiOBoaRdp8LALGeu6XU/Ps3QuQglDP1d/j2Pk7b6LBC/GetA3LSVlByO99MrFc3jT
Uis+PeiceQfBqswyMYaYWrX9+vHVJsNazWa7vgo86RZxlnp6gK0DJSxG2WRTJA6qj9PqQ17/pHTg
a8vlHOU1FR/z0d/S78s/Y0WKoF2NDM7xUBuL7ENDMo/EpoFlV5vbu8xWX/WnmzCinpzUinrX1wmx
LfIoCSHQqDIEtYglSciL1cZWVfvgs4nBzZJh/W0BhnktZFm+owCy7bfpo/uElWTm5UNk7cz381+l
gi6epiEIzeWmvwBttAqEMoyVUzVxVswVbZUmh9D+qz3Zxe9IWOicntxqpvRf/DDILEUKA8i6xnfR
I1/YRKOvRASWu3zku6Vs5rK3UEKW6JWqp+HxZUIxkrZd7IM163eAz0auPze6P4+bG3tvh1wHkqNN
jv6uU3BCThTKIkVlWiMRPZOZkIwk53t39kWSiW1thcYkI6pIne8ffsvVWB3cWQ0FFXDPN8NuUhnJ
qmQ747i2J6Pdn0Hc7G6+BcjdYqrxU785Lkr9QVpE0MVHZsN4+Hh3/jmhzd1267hft4g6T5x0NIam
nn+qpLBLQyLVwKHb4dZ9vNe5D3GKSUzmJLakg5Ef02oB2Hs2UfKoIYZTf8CA1O1lsF83Ti+Fd+lg
eiiRJl67jy1VszhrPM8RyTHb6YZzCU/9lwoR6PoLlvkiE5mPjSuHynrLtDZcoC0tI62MpQVB3Bx0
A71TzYKRdnq7TCqOaL/80BWK11OcMO0KgUTX9nOv5RUzNeaoPPO9D2kD70LC/HRV908spk8ZoJoR
ujIIBwOD0o9Y8RCacFsrFm/6QcokHmFQOWR5zn5ag4+eptWfeG7sPH8Ki3jHrl9PeRp6G0RnLGzS
uwHDlw6RzMYUMTOf0Ps7hanmk1t/2u3GGRGr0QV/AeZ8EukwsyiRFV3M7C0uRTQQZvXUNYU0d/fK
Wm4tnIZYfQoviEolxOKw5t2vHcZaQNC3brW9iLcW/l9Tn+YeKb1tCZdJHQWRGWvV24cV17ckEnAa
JzZTqSSGwv9Dlbgr51mSWWy+KboqJgNFyGOOWqBqaz44ILENZmEKuF2mCTyNJNeHHIzKUhTh69yQ
pOo5e9bW+n7Egzgd6NWoJDEUJoaf2j9L02N/nhfelN+Qbf8sIwihwkCU8b4z/ysbxHTLnBqbY4fy
jOvkwImizji5zY9maSxKygYvhMwc6YobrybVPqEgcIuaQ750PPziI9B8Mn7aA+xQWvbj0rFF7HlR
Ts3seqHAO1/zN0yrOj3BU0cxUwjK5kAcv5v/MRnHTQrOnanRqL8jaEs9uRv6f9pvmjaNuGC+IObe
JWsTMoRGUEuRiL1gLvmEdLTPl6CLfox0yfA2m1N+gRY/cK9sIJ4Qy1vY2a6zLcmxuOAvitYw2G3Q
+cfmOWXe7YjYP0ZC7nEVj4GIT1ZzXoaFaCHBdBzTiURNp8u5hmzqSIU3MwfTUa1Vpy9t3N3VFFJ8
YKvowQ/qUVVvhCYV480Rg2xt4YC3tEfvW/ZhNPMiXi4wEPt+lvDAkb2aeti0R1/ZdyU2wSf+6qi7
jG20ExhSOxNnt87xFKWUN1Sc/z+6BrLKP5toGN6PpwxOpBf4P10N4Da6n/rYatWxrYOt7UINcVcC
/PE2SrIQ+JJ1NN4lsEdjjOJiHhE2Xa2k/ket/+mQit1/Gtr/RP0wuLvCqXx4N0q9czsFOy9ppDw/
OKn+0uTLtZ3LxhR1C3a83LRpiBFH9TMSQ0nfnSTlI1IFxr3KqIkYO5QaTpXH/iMmSIbUv1j3+mRj
TxX/wfTzJ1e3jq3XSHeIrolFyJwPL9ZKD7VGsZSRG5knElMJFh7bj6ylK2QvJKOCCPI2ug+ilmQy
tg3yzN5AtqioNs3ss7G+kFTf70S2EGOEK+tgtxk9kQz16vf9e7wrTfIrbhpGk6Cn7FGk/ARK0NAI
LoJpwWw18MFLy9u0AsFuh0vfG2MzIklcIcdH1G6xsSppQ8W71EIZMdV2R2XHG1ZezzCLP24OFaFU
8NNA6zB/XuvggbmELArDXWKAJqjfMtl3P5ZC/jBelUhn05UEKpyNHXstliTYn4tYDLVxA3Jvk2Xk
5UpZB0rq0ayuUjg9lOIMhNiroOTdhDvzXUmRfHFvPYBhniRpHHi52DtMD2hquQ1ru6o08DamjbB3
sIbeqC1ovXZ8CLmK3iF1TWL/02HBTMclrYoysEEnCOG/HomInys4GY1EBODLfV/zJoNZ8EEMPvW2
bEtTHCjQkHnePvWqiIcjqFoWcFG2RWvCSP10R1YGm+YiqB4Szk0JpSF7jzlgQbc0ZFd+GRRdegIN
hXfHxfk/8X7LA3w+hsfL0DMgs92kl3WgyXL3ZwAQrQh7O/eiVNyTqB1fPU43lBuAo6xNKg5xK3sT
VVESLqhUgGboG9NdYYHoc36UQ3/6BksoxgAKd4ttZpLcMg3mkszyDaijYDMwfcUdx3pQelrt0Koz
80KVna8AXZ517e9sa4FB0yidVCElCe3ECi8pS8c/D1UHSUnuyrVyczKAu6UV5Xqz2RQ5+GJS9VBt
0WKJvNUo64EC72xnMzGce2mWyVEcqbBl/NEOt7nB5lB4+K7J22F9VaocYk+SYBD0NftNNQP8DVkg
SyBYYguOgsHkeheqLONRpgTbQ7brGwIJTzfvRMpU4gW5MAlPWRjWJScYw9yQVYtoiNZ/JTG+MQRf
M5c2r9GyP8DWYm2/W9ss47OAT2dM5YjKWi5f0AsZleTX+ibD5v4CM+CSwHmstBhKdr1z8r7PPXGe
kogzoxUxSHCjbxdDsUIwAq+9qOVHh16Uz57jvRumZyznqp2eTyOmmiNkfanndmXBoQV2Pzlbgqhb
K4qIWF0xqrFAkl4rumF0kgzIRg2ZvfY/a407hvgTd4BKU/twRCZcCjr0k4z3YDZOgCPs2g6jT3u7
LXYK+XXDn1XKNPT7LAldKNK44sopz6f6zfDO/Gq47YZa8COquKxNb6h0VdDIWez5+ueEQawaO1+Q
p9CKFyjskn7ZqGsU4SFeWoMnqikta2aLud51sgQaf1ijUU01DmJWJhS9qtUUyiVMuG9vZYQjG4KR
9s0jBif5s9vN4KGIcRbxcKXRD8xdwyxk1H2/n8lxWiDE9lMROMnfLxuj3ZlzWm74JBMUf6nZlVw3
JQ66w4UAu67NSLIemHtAJvJ+5kIa9P6vg6P9wxW3nMffi0e/QTtvRf3MQJ2qLHN6QRLFx8fqeUCl
G62M9K6cUUjZNB8AToTR+9oeqkfcoTu4LGpyylkYmc2uIazulhHISufBhEHg3AeXIA+FAoMM7MEU
7z4VItis8yu+1/3EeeM5uYYcE/XNhVWOgAFGsenaApbWFuRDMduVMWI7xXviBHLbxLkcCsdTwlmQ
1xwu9LWO2Dwo4jdBILf67jBxfyLc5ogEqFru654Sh1OlZg7XTg2XSCIxpOxtibxARKvRUYWlWMcR
cpApp7urbNiVHnLVE+wIoW1qQj+nXzdwzJmMWEn4chzzFToXy7M9sSD2aVtN1b7b7MqoeDGGnrn6
U/XlJjcugevDpTY7+AfL0RjLecahcfLyuwN/9YIJo8yyJJeYQ6LjCIhC5GD7IuTlZdI70VzpJiNb
0C4Ikyu6iCwowwHEH2UMZc1EIGamhXQ7nmLHNG6WDfU4Nzmzms5WX9/f3XtCFVFYugKGlZC6G807
2Bsdq2XyZxN5bo47iazsY9qpl+eoGvGMUhv7xKGJA7IR0zehlFZIggv+AhFM30tVAiAup/vo/H1m
hkTk+l3vJCbTr7WTz7aKSlR2thz7NqdikNRYXI4bUzQI+OB/DR1ORYmt5PaTmQKWHgOnj/DB65K9
wwcrsEP3p9X9AGOccrM0jU1BW6Xl4fO2JOpiFK8sOqd3iHP7K7RTfKuzeaMdiusqhgflTRyTBli2
Fm/zczFnNt44mMv7lGgnm+5S051Qp45woypKIJwd2JoTMpN2g/qgBQLkiiCh8ysHoB3DEbsgsemn
1Lcsz1T9VGVp4s98wicsMACUrr8knQb9ASEO/A1Ctgz6dZYoNM9sA7AAGWRShP+xUIEW45qGlDbK
sHheB5eoRbpEVh4Qy65XDF5aOyjBnKm7gCe3IYjbBJkTEFlqXiqzAy2l0XhtYyMgLFurpjX8ZHfN
VpqIJi9ZjFLs5g6WSjKKTp73A/kco7/M+AX5mvwcjacoyz6wsoZrUDUGaqF/i6+oJIuiZWzvBekb
morLLQJolEinF+Mocssx+Hda7n9YS8xGsUMPeAkJrM7Q8D1FDytp6sjcKtnQBb5M9+5WFYdFo1fR
7myPxU0cLQ+VRrETie4HwssTR2Y2Qg3IC9UZfgOiabsz+mjZP2hbbybhCRUr5qAk9hoiloI5YIIQ
0zZa3nUBdM+hAluEfYqTsHPvbMtrzIeiNTy9yEZqXMcg76xmeO1e46L/mQrkl/hV5zi0V5N8sG8u
HhIN36+iz77rILbgUl3zm3508gbLM0AbErwKOd7q84G26gDwjXGQBuJuQfBuQ33TuxjEJqIipQcq
13wM9jZNKlVdPww7fxLY4U/8Tip133z7nDt4tTEHvDJYrELbtLS59B+LoYJRYxzcV3WvJp9Xn0rG
liHac4iAjqIQh6s+H2O/HyPiCCPvZ6sJRCesr/dHuRvhSDptUiY/8JTKwjZflxX+0bs+wO1EtiKR
KoVTOWFqrYDStzJo75dDAtMagqiFkC6Hhu9m8s4uPouoIfxGym4nG6YDdzWjzxU4PtuUf1cM8VMp
WIuyWlsctiwkmLSoXIQsncPurVF+abEUsjZhNr941Sdc3dAgWY9gO4GUDhl5pja4GfJFtCM6+pLH
LjAevVRMYlOtMjPGY65KM/GHktJr9177TSOxQgYUQXCtHUsEqvFLj0gjmHxik9YjMWu9t8mAqkgL
DvTHXg/3/uajkcTkT/lbJlCqy2Xo6zLF0somXPzzgW21VOG7r4ZvccVdGctkvY5rVUtGieHlGDuQ
kAX3Hqy8I5zOFOS/iN1D//wo0EbhmUQtzEqbnfKykTU60COBr2gh0KOwy9EbgbX2H98yuBPVc9tf
JHM6YOtHTQz92oWWpn5G8a1gCjk1fGxbk6emkmwXSVx9CHTpVPdurNioc6OwOkulsRf35umK6/TG
2fU3e9FIfGgcc2BOLMaMoSE9LO2qUItvMUtb8c+IBzpLtWIMKYZAUjmJ6eUNCUOGlV0twrhcRN6s
qGRels6Tct0HOTsZ/HoLgoyAQqZBL6cSOAWwUyVfvb31cMYL2NKsxksY0cXb/xvzyH/UjExQudCm
CT9buz7AWosxTlbJBIgZQam3uYNO/r1inDrMGXBKRlVJ6XBazauYzqMKChlPW78r/X1V7CS7lkCB
xo+gzwdU3DEeMN7shq9gtka0ritM91w0tbkm8EgeHY52o9F9XEPYtUlM3tKV+clunOeljIbQLGOa
C/L7Jf9m3mhP0UpuPpMW6s6+H+kGo0ZM/ETxNyQyJt6006rGhRVYI+SrgqimypuLNHo6pIJEVshu
c/us+yPbu1Cu62S9dmarOLxB/7uo801q+Y5LeuKlrI/bAdmST0/qNTgKnkxOePj30BctK0yvNdm7
qLI7oVQssuMj/1Xy3OG1B2VlZEo/kpu+piDoIKVs8iHx9tbYtdHVNkBNcychHkDFBa2XHZZHykXI
d2mBaFX6sN7MfUm3LadXThBAyzvKfUZCjog3p5fDLypx5utvQfvGO3QLNc82g8VTUD1zujlmlzSs
vxlwgTSEhsYBhZpB83MSbUlbNBdXB8DItQKPnWERoaCV6tVZM9lHiRnF/OTyxoTVq+eUjM6dGzPB
+1QrF/fasdeH7EF/ljoZxg4eFjYcIwvmb3Xr4/TuHTS37pQwp8NwIbvoNw4wkHtWyrQKO5PCy2bK
V17ApKR5v4WCmjMLyEYCVG4EAgeoELkI5/BC9YOixlMcZ63z52V0UBxgVy9lqRJZ14D8uSCJ1KSX
s8QEsHebzvnO84jNFlHMwR+wAdgoPk+0fOU5+2TUe4pL9IufCZPXXDT3gn/an58q/3k1scyInKth
M4Lc3VGEYjw0p0foS8lrfwmEnmkzJNHEg7k++4UFChfUUAWPCpFhi7FEG2i3ZQ2AUeOYZexPxBH3
GubX9eyyPjqxdPFxGHUfzT+T8RWZXPGR+zQQb6PU0EiGC3z7g5ehdOMhdPyii+M/GsqhjqZg26yl
CCmLrIIpRbQFxR5H3JQpvbQw6wDDJyP7gtFDroyeoCl4QQkJuGj8j0YSA1xxgYucgVoAvVMUs8xp
rpUQJqsz1TeOmqp59+nkMihwYt4GAAb22+I8WVb6PkUqs5F2hDHmI8vb4I4CeC3zHpxOq8AtBtAa
+4skncoOqFAIaSladpPSupTDR5lFjZPxalVJLEo7ZDWEk6zpxu1xc6Bn+tz1Sy/Cue2VkbV/ud+R
HoJawMGRB0aLmkmtDnmphSKlrqZkAaWCrlWCwLiTLRN+kV63egY0uHDXOcmtVUpky+ixhFQzrXKp
zmvz6kANsS8Ts5sEfgbfka70nf8HTd3diGH+NZd9rD9j1gOFwsa8S+HtyjZ+9av81aUPQZCBVt7d
0GbUeJ+eYJgBPWKzGFy12sEwYHeDbaxLoXbaH3wVJNaXIyeUCzOhM4PEfuVG9hReijfnlo+49h/K
Cefl3WO3rRHjnnK2sDvYlfsRMtF6gd4bJcKaZ4qeFla0Dbv6fQyQ727QgD6hlFUSL3biW/Br6VzI
UJMbKoltQsWPWbNe0GRO25EQtyz42+q7eNL0FK4zuSCroEf2m814crO1o//zo5OSBc5QiOeqsDiL
WBgUwQR2Ml42gGRxRruNaj/f7qOnKJuCTYt3EfO1CnL/5fBPWzZfqLd/ZhNoPAUVsjATeY1CRlTU
BylriwvS84lRz5iHbM5SvOsqWtMDmDbn/JKKN7l0EmvW6nsVgM7q2+UKIgqVuiALFmH8xx3lQDW6
NFhnpFc2jdi9IaEm4EY8xe5ftENsUf7ggf8596YZvQ759Ty/SvRgSYmhPKTJ9Qw+8FXMhd4U3Nrl
YU7WTzfcsMWRDgVfx7uCf43fpe9x+9PZ8EMiSa8BSsZekXDLxLShgPRjceswIAFy03ApU/2ng2Qz
f8HzBTXxyP/09tEF7u54Vu54cIK7KtjGZ9J5iniGhGg9lW0RxQoU276rR+keSp2Ra+UUgD84y5Do
CtUffHdetumii0CxysZc+YTB0UFqxQRiAI7JgIJIVanzvjX4z2Hgqg88SCYfmg3Me8P+EQkWxXCY
GYMUF9IYlBwmpt7ENigPYpBO6FZqMQourcdz2FoU/J7izEN68F11cd/hujIodjTXCHK5JePEoWRR
PGqQeZvIGNIec3jh6RPetyr47GBL/C7aZiWMp1tGicgJl1KGGMmlt5EB3DehzAjelqSkSmK9Xqia
rGzwNbuoeetbuN8Kr3Q/kE3IcyHthgkK9VUvVRsPDWQFZrCmxN+Lj+Jde0+NTlfH9r3J41bfZFYR
zX9WPLQpAcy40vDKNitPZjaMdrcEoS2tXVLaXiruCFgADVkh1ZEbJxdOEZwffTdQECeqrJTRqYBS
VMr/3hCEoAuWsn8lbJ4/i6Hyg4XxgbTyEJDmEt9JOKsob1qnoY7lkeqP5v5ZqDsyRyfFlL53BdqX
fVEP5DgSF0UVBDxvmH2O8hnWMl3O0X30mOdr50k4UE8knD2+xbA6hKFhB26hzvd+1QygDeiq4BJ6
mFiiV+iEdg8zRIciclniDCz82x92oJyuLOPcnTCaUSen246Y5EVMjeMCgDI57L3/3dkc20VytLcx
8hbPX3L4f78Qk6cQJuQ8i2NIl0wPzPKXhzP19ohN247HyY5+ip8LAZOy2PfWySKVHt3K1/BBCoTO
KyvdjonWkjewo3lXQ39a8i549EjtlZRZsGE7JQ+P5OGWtAZnxsd0HxsWNP7kMx/VT8vzZpVk1uMg
YQ7MfLu5ZXIC3W0guDPluAphfRQPNxU+UmPhZpW698FkDxymEJngTwjLP5d4qcmDxy1KZWjqaW7E
07LmKECSriYBSBUm8LlH5yJupyrco1nbNH8YzZS/Kof8+Nt6+JLrmfevjIGfdH2DYSCce9yxOxX0
M8J5Fe5IIE0/bqSQlvEiV6EZasu0RyzMY/+IWjcQnu3LdImmpZajOjHmSlQZLv8eczvdpoJfzD71
bgfmWH41fw2ly2WYWDITCLb+lQxtPq72w2ZRD6+qwVkCh9HgYI1fyXr+HHyfErw2hQKjFNutB5b1
Ux5opq7VIoy0F3R4xl94rkE1I0bIWuOlA6DnC880RfTo6g2LgmPEbJi6jPpvSV2VKviTJ3NDcI0j
cxPK2iEiXLL0j6yyHKQ0Svq/cIodiEpI3rYexZa5V4yk0DE210bl75ACL1PeOAfsKeRm4lc+FHjM
SDRHUHBO6h35TMLsuhmMida/+r6ghFau4RzOoSG7cubYp6vdoiV6f/XfpLGfOENYPrTsGKea905R
g1e4G0oiVni8ASo7RqHVkfcHmuy+nuLILVsVSc+qmJDf5tP+KYe31pa46SzOou44IGy6DFnq6wlc
ax0AMULOxK2kpQ3KNtJ1nM3M3OSX36fZecylFMsSY8pv6I9ywJJjnkzRivwwicMa2V0ZL5xlTJGp
7Cv9IJyIwCuKWX3VlsuZPjFoWxHAMcwTGRzMvFqvwZtK7Hrmc6qP2mZEjSXC5Qdci5Z2Vj5yk6kp
JDebWA6b7FP8+R8agwJXqiOcXIVwhCH+KU6ootM7LKoKblzo7qKKc47BJ2JS1KZA8hMfcuiQ4GlS
/R0ejCv2Ih4GnwCrn/bWLrehOWsdk1otYJKrnzmJ1YOzjpLtpRlu17dlnfjK/fa8oWwJkufxnA8m
Om2BBM+hlefKns5y6Gg4jbVcdu2I9dCPWaSan6W/IkKFdQUDm3xIQAKjMXcQdR0I+9+hPBdkySVL
rOsjfnKua426XCr4BytDi3BJJV0NJ3g34dIVOM+1q5DxQQuSciUyuqm4CviNnOulGDZjuXmckMjB
242+t5KEt98a64RMdesvkfifQ4G9whjr3jIHQcx6AAvTx+LA21MgB+pYK8e4ke2xhTpwAWQ39Mk7
wft5OD63Vp++EKjQ8YwWTRkTdIcZVdF25Rbm5O97xN96O3sgGW7SGgo21ZOulpweeZcDAQL16rGb
se68Ts4FdpIU30+GAiCs12/jzEAQXN6SHrPEye+qjWqk7O7t9dlHbPULCq20tq1XZS7tO9FODfxh
WfLAfJRFezpddVacivPrG5rPN7YLshsqdNCZzIKZCVf6ayO2qfVIG11+lim83buxrGxQOjGe5JvO
eTvWJvCk189o012ocdzjAiF4BY9MvyXyOepHIiJaa+3fGTUd2R02uDZuKjVJE222q3UCa4lHutvi
pv3sdi7rQSv40rw5qsezRCKVVUoxtLam4nYCzBY+bYB0VZbazV1HkTUZgQ6uBRqVXRDUku0z4OvB
okpLcKpIDidx+VpbYleJAKET3rva8W3POYJUuSgKRmtCHkIjyK7PLEbC9YtZ0D/Batwj/D3onacj
mSiS5oA0xxRDkLNWW/neGmUV2NKYhv+M43VOXi0ErSVQZcVhk9fMEg8IDoaiAWPwA9HpFlBfkikP
qRRql0z+F3/OP7+Sph557IXRP3I3mDTJjBZ0W+cgu9s/oXbZVFCIIZV9EkwlZ0gG1ZkyWFyf+Q/N
/q6MIa5oOhvEpPshaxSZokIH5l0/VMbLsXXrvhJsyb45K97VmsvYQTPFmbBy75khA9MleGuWIbQC
TSRcVQ+ZfviUVbh5iwTjuwI+DhZuYgrodeYH1NIEPs6Ac0LjUro71XHzS/brPIHWfCd+6tcY/hva
XdKUVfl6fNcTAngyr3cJb0uD1N6aifEDDC49/7qfDpONvFLUHZ7QoNsGBuUbSbcaWJS3jyveDJ+w
UfF/UMXRdROWV0tQxnxkpLJzm/jfK3Qi7VfMjGS772jsHoKfD3uRe+aSoIsZuSNWE+j9qlhJcwbR
SgZhoxrb1K9j6k4zcRCRvPsXTlvTmG6tOlLtPYWqtmWWw1+QGP6TMQ9s+QQdysYyF+P7HouUL5zL
dAALgikO5iEqcn7cUCh7OKUwKBxdVYZH2b+7rqYCWJrQey2d+lsWMYgnO9Z9PKGlmQttxjseGwRh
Qjhq7Dw4EqnUKNq/OfSgL16rm2IACvMPZjv9SrONctF9ADj5U277IZ5iTWMU9YD/eMD6T7AksqHc
7/gzf8r6/J1e4gisgp7kDayWUTL7Hu/8zwSWnbtS5Bve2UFb/wVBzffmEQhVHBz6hPXREBjLqTs1
KDtHKIdp3sGZEBeiz2Dvc9CPbWc7EiQDE5T0VJIZdkVDX1rTL2hIvx8lzLd2e3P5EhUpZdRF/XsU
4KJ4eliX8DIxYudr5vLSqbL/AonHfG1OV2/7NvdRfF4hsKOitmwHNMJXP6L5mRaQDwOd350On3LV
kmR3Xd8b+s5UMuy4nd4+SiuaVNDplW9PEIL2or+dhHICSws4ZEIJvszVRcJ5lCi6GhWYJxllAt1I
YKoJTFjaFXuk2boF0fpKKIhDmGBHvIkT535D91F6yCo3zyAaTHKy9cYuJFYcAEEa95IzAFZAlmMs
02rcyAKZfCvujSN6mqd0Mw42pV6BLNrg9rl00pcJ+xEr4VYArBrn1T4Z86CY8rm9JBeuQz0zDoau
vn1EO+FNWichZ42saJGXTLUwAMobvxcxnZ7rOX5JwRshTu7dChDzPxRx9VhEpJlVsKHmwsd/dLLC
ABvWHU8GQHJEFbU1WSHViQ4m7Al6FruPEBaqwBGqDczjMuuB+S2PERvnTokYnVxI6u3PFkztD6NP
QvaiPe17OMIcpRsFvGWXo9mz6V33M0OBrlMBgfxyuZYg+dbWlq1exr0Xm+knyxG3MZ5dQn0zxi5A
CR/BLUJWywWcqyw92c413LzOO195LnAmK6+ymMrgtcO/98KgUEWulYyg9k8Ic9ARnoYCNx/4eKYT
VrQBeOyyXCcU6T+lMRNmWDS80EvZkXRBm95ktz+1lBPi/OKoavI0Ixpjz42k07JZxuIKlYoz5+Dw
pbc/cZo39TjT5wE1O+AHZ0r58jprW+DcleZttPcbxV+5LizMaD5teV2rukQOMwS4lUso8bke6OtP
jh/ZDVq7kjlKUD5NS7JuLwGkTfdZBdUV1SiFjajJlBizngM5Xt+9d7hWNVERkrNWLTK5StXlo515
Po21GXEvyOex8tg/UgMngdCOUhzCk/2E366pkvNyF7C2WIzu9drxM0pDCA59vXsS3gdXfM6DTA+Y
V+TLuKcIr80wwUj0s7TRLT+kxuSy5FOWwlHYovC/7WdwfnaN0cLUJKKD7PxKHbuqnwc15oSlgdhx
eQ9npYycS9grc7L9eThY5fwAAZ1GCfuC//67xCBfaPc7MTkvhv2O03SUQ3HRQwGbHqf6GRMHeZgv
t3WcSsrd5lMu7TXA7k26EfFzVDyIsEPHjWfYWsyeX37ea3c58XxBoLi2/l6QEiBXKqEfLpjQC6dL
9kwy/zHH4F2w3DSHfbkLqx+hektD8gk55TYoHj8bLMbwR1WSiX58cOYvR/Ifwq4+IzjeOAOj7L35
BiCTSobvrCOO5F+KRtNkugcpUIQYEKj/1A+ZLplWyfHJQY0aDI6bG2hpCU/PJHuSZasXIxQ1Z7IX
G1z9prEgL40DqykJSwwFFVyMuJONzQcx1LkFouAh93kcLhhsGkokWu7abcZ8LM8563dVEXLG3ImF
YlT2ae+vs1S2VuBk8LSaX6dFt2x4tvVL98ZJDzIWOsBjxl+X/XzSJB+pqijGI2jzYQo/Z6FhcNby
rt5h8Cyid4zVnQia2iS7MwhpcO1XAcZVR7crBMBQ8byHNGEz9nEvnz2241qLgpHYDYObolo16nVc
CBIc/AfXbl745cr7BQ8kMH9URPOjXICKTGG49C/F5rVu6bYlL2eGQ6RuiMkHsWSNPcKxlCKl1RWj
PgPN7erVzZzur4HnkcMoB5Ut0+XQHHBh8iFpS403rVlGf4ZPZTqChe8Xrcos8lk7/d2CsAH4OroO
brgjNiP1QpCkH/nX5avjuzKH1xI/boOy+iY38Rxy5l44G27nyGP3KWldMXNz+8qAr8CXrnrSF8zd
k1nqS6sLNQA2s9d+ubyxCO8Oxe589smDxT0DVTBTa4gv1EOQOfR46+RzqDQknkJc0b66HVFTxMxy
YxiatJhUXa7pd6o+nw5IPKkAzV2T8AVAvQBBRE1tDbQY26U4jUscdldfQ4XyNy6m6D0TPkjOYA13
uguvoPN+xbcMHAwujLsXBCJ0ypqQJ8PLlp4v7BC/fW5F4Db6z0bPPZdBYq3sPbfzlY7txqIzU5fk
gZKPevQHcS3Ug7Wqw1tDiRMboxP+7kpJFTdwY6VedGPWIZB3+/65go6Ny2X0+ajEv5PDDsdDcq6/
xvs7DrF3wiBzozkBsPTrXxt8EzY6uym03Q5lLlMsiAwvt/7Lg0udkXDmCjqyjX4quwp6UTH52de9
xEPL7MpDleoNv4hbnb6FCLVq7Dwx95k43wcafbOXs0WmjdaEWS85CDdYuJvj1TRcfZOSyGMurKMK
WZ034Z26G4ur643khmKyXO7pFATUukUiNQC7klgvlwUGMi2IAek4Zl2afxw5ui3jDNEM2UHE7pH+
uO88D4lEqs1SqX7Gl4QK1XphGaYe6DXEJCbPGCsPwpjQaOOC0CWGy9VZseR+L1BVD8F+U76hZUPp
uVQGdT8Htgr8wzGqrdjnDnnMizmDdfrp6YcsU3ej+rnNczHC7MpYyfku/Pv3P7UteeHWqK7bzn++
2E9B9MsOryAnYpjOsVFCklV5XJCZ7E5XZs6MB0kCw1FsPCobTTeQfE7KEatY4VYf4Ba7nw8BZ+a3
wknt2PrUlopXzbfhdQg7h6OOf6b7GSgXx91+h4TWsiH3zsvHSMN1slKL8892fSh14idSsHUWDWrs
SZz0NWyP/AiN1oKGmXsjyFP8PKI4cq9+lWxEKn31PYBUuTObJosS4bApJ6THevub3i872qrEo2G/
Qq/F4yQ5bewxOkZlONbm6CDlTNhmpYIA1jQqiwJxqRoZpleHJPedGaHGZa5uxQp93E/xOQCUG1w1
svbZ7f81EDkh2qaOL6pdTYTEaCvwAn+gD9n7DOsYJ3mqABmXyjSG6GANM8bpHe1Sxzv5EqiQcTUo
qxLjrEjcFmQ615X4wrxReuKaHGNbBTxW5iZxPTMjkQeYRysgnJLKkA++aYVS4jDoMdySSmeQmOXJ
Bg9dJSvX0vmaZjgIbhilyZNywe6w5xvlws7zNtSUOSPSNVnFN/wqeTomjISs9yrO6hSrGNiJfZZL
Gd3uyhWTTEC599nTWDjtqv0zEF92OLIrjT3A3J7Ww1EERMbKPPFHGag2HWiA2cMAOK7v2PLjpRZJ
GkRv8HxRS02O7nzv8cKXgtlR0s98UHPAvDBDWZsHfCQWnkJN4G8C0l38YanED/VLZp8RHGsyA8rH
CAGTUShvjOx+NGDym5N0eyHLi+tysdU9W+1D6Y/Lz0M2Ns9AHWwQaBs/CCyYECpTSvDFJb0ej9gQ
wxc4hFcu1AjGEI7qUP8hn3dm4OaWjTUfxDOWchfCctrmJRSSCWWto/pmfkj1fTkWDgm6fgRCVOpI
Rg/3BuBQ/P0dope62AYBdr8jpOTwnznvM4Ak3Ljg4NPdQVlRJYYme9lBH3qB7Pny0elwWxJDsfr5
6UJt9xKWDzpwDp9SCxAR/Lt2rdtnM3x4cqsmeudj2RbaKOyNByYNtre6Me1v4RQPbwWM+uysaDML
f2YQjZgTiiqSO4QVGxmteDDzre0qaNA9shZ9BhzFkfIbDzUv3FAJSXxFIpCpdDgWc9QZxvOAOkU3
hSsyc33SWhygTqmbqs22QKRCBWtGRKSGktjswVZY78SXddGfQ2w3grBgS3tlLpqAg7uQ73TMiUph
MgXK9BS8Y6u9Xu1GkUZBJNnaA0lztBZ6wZ0DvdTbaIDIrcbPekRxgrX/oIQ3d/n4tCWYB+qq0TgK
pX/Qu4ozvFLF7+1wvwdzZyFSM9RUjV2T/roRPvIOJ8KAdqd9IXsw+nkUifcOX8EYtUAgmUkt4b2P
CipY+B8rjaL2f4/QdFCkR+Y7cV+AT8Ez0qBQ85Wgp9hkUFV5Cngm+K9+t36h7JfeO8IP7kh2pJmI
WM4tdNmbSxnRhvub3oj0/FkFiCOvOFlnijxkg2F7hDtqvav9aYBVCLQo6Q6WocXbdX2WVTBKJYG3
7cZq5IwgbkW+N3isiH8JxGPcszw3LgxObQHfJ/YdzhaLAoi8AP7WQY8SChCLSYzIU79ZC1kBv2WG
rUfSZvTXRnLAa5D9NKgwkHYyj3ykBaUXq3JaYbyCvp/6Ysip5jbFM47md4nulskuyIX4Qao06HLH
RBp2UJnv4MNdKdPMXoen45msh2mdEN5nuPVOd7N7gqj2LrkYkcTerHg+IjjXNdPTesNi1T6WA0Y6
mC17zSAMiuuM9ncghX/exwUUA59l63AS6zZZUT20upj6ICu8l/GKlyqPtlT73Scu1CS5r2cA1LMo
IXr5DcA3HqVfGgxjI5BhjEGuGYZg/EIJv8o1zdc3iXKhFgQFkDxnRtbzbIpIjVWOuskxoPPOXuVW
YCd5SV08VcETmWRfS572L/yfPFFmK9biWbuCu9RQ7PYGua/YL0kHE/Os+2VVCWf5jf48B/0y9CtO
wyEAAp2qS8ACbRRVAYAsvDoLsL7Pw0agOV0/kGFHPmrjYwjZkoW0vdZnjrosLb/UW6oY4WcrGyg1
VkQKplkKvX/gPfkJi8ZX6mbZOX+ZCQjxX2wA+KCHDGL4n+PNjDLTQdYBFvn5RqV5AfzvgLoVBYSh
rMyC9dOoat1pXaeRV3OmnfL2YDpVqsHbDZQtMaO419+4+2HveSuJqgtB+AgauAzwvetOnrKpOfkI
miv4KTqmUKA0HUWDnFN8uJhSobDZd9DD/1IZ6KcEubsGGmXAApKAz/XO6Of35+6yqKiA1Qbim42f
CE8A97+BmGa42dIQk2pVvbwwlBtnE/FgmdxZb+feTqJnGwifMUd6DpBsdKHibqX/SMvQYwPSokuW
rOxp2swTGXcuyvDEozhUjXIk1eKpWE1swXw1KCD6K/jN7OGh6uRqrKDzab8ASf/xPsQSPbmqWpfx
zb/BLobZh75wcBnLUFLLA2ANq0DFOCCdXpmQkWD5tPUQrkuBSYts+U/Sye4jFzDbCI8wtm2nrt3g
ruX2t5P0lDyx9ngMlSWRQFhz9IKPGOZzk8Ts8gVgHybn/h8dU5e0Ts2hLeMGTEiNJ4g/arbwlw3Q
pW8RIz2+qeolRfNWOPdKEox6Im1i/rnBjph/+U1EoH4n5dI9DhPsO7LFOzE4KUEi2k3TI6xgF/bh
GTUM+Yld0jhfoNgeW3lr1gA5YWrcCoHvA4M5mHjL3Rn1rHp/0bJBiPYGJzBqkxVu0TAAViTXb3sa
40jlRZL/VRy8hRiwoyOFFRcxjqoK5dW+5PZDQUiFV53KCcl2DIQfBsmWAtcgrA86M9qJHdJQ+Blg
pHGoZ2uP/Ic+gutIRkKrqlWigtjxgiGKnzZaQlUsI93QxuHxcNKhM6aXmbdbrF1O1UT9TRCCnuE1
MaNSQ2/5h6sZeAVqFtKbH1bGwOaQ0wBJbhgT5df7qOesQgHhBcfVcdbM6Bsh5191Guz1XmYjEJh1
zDh4U3UX7m2HJBsi0cXua1HJJnG+ab8n8bpDZO9C6PvBqCbufn15QYQd0w00YIMsSZnuIFhNoUaZ
/2G0wPPlWyv/9dTEeiCv800GYfg1c1T0izvPPr4uMmkqM8+4kkrp3vrH55ZSH78WC1aw8KOytSb9
R8OZC5/DZFNLO3QXCxsW7dyLkRd2Rfw9cmBw63CXxNl8HM1wXA0Zud5WsyewopZDdSWRT6hvY+8L
34ERREfm3Uz4dXszv02AnXE3syd9Ogey8PwOm20hFUAeRoq9Uv7I4nZ18lofNBBl43c1l22dNbQc
ak4q6wDDBi/4N9RYrGLZauaCj22S5evyvoICYbwQQQ8m+/mUZALLzuc8hgNMvT1aZm71ZjY4UJSD
+XFpriO9P+nLPJi/z+mqYB4yfxXezB4PjKWJ/7Sb+gTQ2BuR53cxk5BtYk2bdQvq5spM0sGzkld8
xEXFLlQz7duBvmxTCnCtupcQ2XCCW6XrG0IDkqP8TJL9Rwi8PUelsPEtsSmcwnc5J6fQZMlJ8nUb
N2DuGsf6w9EvSjiKVHbYonnHvgy7LOHquUDq7PIB5jOcgcceYfy3joHGIU8hBxlbVl4NPmRvXSmA
IKLz80cROzW2aA3dT//QCZ6+YJq6Yh7QD2mUr1kXYuFyNo6nJ+GNIblRucDrJV/jhQAmuhKIW3sO
Cr/tgxmQMmLEqZ/hU1xMI72sCgZBJXFtOhevcQSNgV+Nn27T0Q0TNk/m3gA6r+V9o1vdopTd464c
m2Fdc+3Ywl5w3P+GUzVo20b9d3ux5rQmI/fDT69yKT6hPLQaY69mrJW5ahwthKHqQz7bvKNXkyZZ
fEIHfFb2C8fMOaRK/qk2/rx1oOA2WqJkGzsWrPcN2dXZ9vzMGU3OZLoKUfQ8MQXrvAeQOC+ZfwDp
+tXhZBWiOY9ychzHzkHN+qC7gAohhwcVpTk9ylgISPn305JyzAEGelqbSaHHdKicEoXOLbmjrBG3
lPpDII5wj1JKZ2hlV7D+zAvHJSoR/9vedYcqlsH5JqemNK8Zux9+Zzc6ysefigFmmorTSVltjOFt
hn1dWS/3sK0kKR9VOO3GTsKkAvxyyipKNXI9RmW5E1YIS+EV1fSlGz4bnZkeMU3NjfkCZXsSa+4I
Ku6lEnFaFtZoJCtOI7emw8sn7HCkmjo5y57D/hlgXhDPG0Me2JvGqgxOaCphi9PfFm9S4xwtLg4/
nl4IdWW9HywDuiHocl0Z00hngfBpQASdZ/c2AWZqsM14JSp9w4/SnD9wu9/BjuZNoTb7qIAe64nX
tyyj9qt/sLVgQn+qJe56dFpt+mbk58wwUrxWyIYnfH2YkLOxXLKDgfXuDand5xZdvBknARri3im6
enWwMm9qHcK75KWA8RaoXdyZSYCNiZ8lWD56N13VLNJYEfPpikXEf+qGTEubC5WnnwKSfzo87kwO
nwkSLtjq87qKTo4vD0WMnuXjBdP0/iI/XWOfusyYj5mCz+RNkwjciNpMHIQIrFzq7uiLIo7aByze
HCNDHyt+O8m96fHxSqDuwotpxcgFt6v238j/3ft69VKxg2EI0O+3H60WsRSOJRcGIOtf/UpX5yMf
S3W8BlWDhgfZnqEKjWt9p36MOxKULASVoMPSv8fLAghp/GundHIQnNnkP8ggGcIOrQ2uM1spP035
qDWHWn2B15w17db9lDvO4v7PjciDRtiUi8SIcR5VzoC1pnWrChUOpbZRg2GMp7TFdSAckIut6/5S
tfDvWAZm7QNKIv5lDbdX36TGgYnTqhoyvNA4ve8peCMGL22e8zcTknDj9jfXy1C5LmL4rJGIqgBM
kYsiu86C7Cebo/r/aqhTyrc1nX4a5B8ntxFoHqnvgI9hlYqzgJgXSVFLsMHPUyk64eGt6WCkXKxa
k2oUUqyGZghtoitYATK/G6evBJwju9kThq3oj62V7VjlceV3dc9VqwRYPmpDtNUUBSFqrLTnPeBX
BTlJLkwDGtKPujwftnE7StGJcMfxuXdpggu2MJpa8rnLGxqIH/oAeH4/9xcTHaW4IvCUIB0hA4lS
lsLDHDTBfQHlFpXl2Mc5XOCyARTF9Gn13qXWzUMbgsRiWLVvVGoP11TAlSBfmtVsVndcRBTyAgiZ
lnburbZzYNld1svrpzG2VsshOZGJwoUQrX7PuLD2PMbTG8axSSYSBaNEXLrmvqexRtjN8ik8XF7y
1yyPUeazntqiEr1VfYXaMCtBRG4Q5n/XrAIRR2KmbuDtC2DmIyrLdsmBNPaJubONiFTt4rZySFzf
10EBSALeSXoiO13l7DaR10TH0Q22ErqpvyWRkHcmZ2In2KcUUNKlKYawEuDzsu1UQUCPW46+Seqc
J1Hlqf5pwzgoLxSw0/Qfu7bDkloSFs4SZy18i0i+zcdjX0pVKaGgY+xyAzHULLXy8rCY5BFeLMfs
6kVraF2/SCfNklmYW2VXwciwDTNk2jvsHKcQE7TwAH30ZP4Rc/deF9eoYy358jYCmXhcdmQBD+j5
6onlNW8qSIJBQpDZrt5NaUt8aaWQ7hoF0YEAmvKVtXhzz3dfd0SGGEruo1VHCcgYB6uIBtJKqowy
IzO3gDlfb5e3al6NvSmRUQCdkI8iB+nEcJqZ8WRTxtQwPwL/0ILsCXEWXcgEMISKRZYKKIcr3B7+
JJ812/DhTJL5Qd75tblcrsP7xyx0VrhrIXoSl2UwXAiktzJYWCBhrgZlGlx4yqeMepUm+uEBHwIC
PjMYiK4zuYZB8s4Ne16lLDgsul8/DEv05qKPyMJQD5LNQjWQX8QAK5a8crGavo4O+eyEJ1PvXyRM
hHYjfp9O274mLpveR009yGxtzATkXUtzgryyayV9hcWCtz6QJ5AnI++WPY7qKEPJyo3TDcrbO8tW
pFu6x3kYjy8pdRb5weM66bgZrXV4d69CVuZlKrE5P1vUjgRBEiru/I+mPeXs/O7x+pDLo/RxEiiC
j8xt1gTk4tuTi0csW0/g4tqsgVr5c8TuTAxE0O02rWb+B6yihaQTdPoPX0EKKqadxRzYqmczOvZz
x9Z4l9HziEJs6nxS9LwTxq64kgezxf24iawVHMdqnIzVDwgfzwl9hVnKS2xXaPJrKRodVFz9e36b
Nfs/mNJtz04hjHUbkB3yFgwn7ryKb2uZVLGRPEe82A0Fw1ZSQkyFa5c3F4UmT1RG1O2n3iddcbDv
U1MUHAxO4dQm8By31PU+94oseBgjJAv2Bd2jjdIWoMoCKNZtqrtXl5o6LnlsjQZPBqFqd80sl5As
XREZeqOVPUFfvQt5Tj1lFccgXeGMq6PNTwYFcUjMXDR5vKwB79skLRi1jjMecsBvxIFtABj5N6FM
AuAnJ6fcH0hJSfFoOuNSyEOuw4E8681t2BISBn39TcDrkSURWzPilAONmiN6O2/7v8cS/HLYqc0a
BrRtKUSjUYR+rkFosmXfkxBBiK0dl4ImdV4V+2m6/P8NLZNm5EGi6E3NxUKg4pVROIq85XF0rgTD
60CGeOsP8GmYyvwWvivvLKNRFd0uhBsLEGjK890PpDLVDLBzA8Unn5PuhVzKDWDqTt8X2004WnNp
0wWRuI66EFoQ14xA2Kuv+6zYgXVc00YuOiPieihEMvrkY8pIhIKl0my3Uaqu73gHcRXs2g00jCT+
PvrhhvXqhEt00lQgrC2mdGGak+9onVq/Kft93ai+KUY1ZoGe2Sprc7G5iDv/6zxJrzvc5sMn6kdh
N6eEzew2ZQ739+xgFXsSJnLbvfoRh34UUcAGpgUFvmrw2xnJ+jUsBR73l7NSxaVL9xJiwvlm4uFF
WXNqx76BikWHfDAGgAJi2UG+d7kMQ5UXAH3LyXclZGK/CGC0ZtrcW0i+tkR/cxLRqNBXbcyp98XT
azghGLdyQWIktcTnnuyteh/jk0HT1gg76YUsQW32Rb+sw/CxJlK75NfhR80EOSTj+gvCMTHdWFsE
oxG8HUQSKZ9mynqMRMJTY4CvQfI2HQaz8TCJeEY3LQ2w25IWibTTAgG5BdjgTz9yAdRKW5smbIe4
LXIC54IW2RMmb8fyc0z170EdPG4P/StmEjxd572AB9KBt+XABjOUsZjn0XKbn2HdFBg4VsrrOM0U
iCKb4fEgCUd2HJkMyUCpLJ0Q0Ndf61/1xccqaoLVvIqtLc1yYbgq/nGZb5SXZYtYLAmQhIzGhdAo
+YGrJhrEkluW5i3PJGeDkDGm2IG5367M45xFjkVxctzLQf0iXi6szzIWQqAPGvvDgHjUyxEeZlbL
j9s2gUIhgjfbjnt5UZVA6kyil7q4/rYAGge33nvc+h128jLO1jvmH2J7TnknVI675loEDxQd4ce2
qnwUYMrlOa4BCsaCRJtMD8bSL6Tvfe8ayt0ERdAG0PO8I4oAnKa1GZ+w3Zhd/8Qx6uswZZFjTV0w
w68SKhPejYzitlEb6HaP/I2gZ7h4oTSGAISVOuUT58JdpTMYYR5wz/KsYFoppOtNbLBBwh/fi5rX
exEiz6d5JVhwlehrhasvqbOpAbW+YDSWhdPbyV0Ih4DEttCGATlFeNtGZ2zWvS6aBNMXV9F5SgVT
hIB91ioKz5IRiorL6/Blsh0WthBS6Zhu11+oHhNDxh4GxeOmkUcMTxcvzgDnqrZadbrX+rKtaMHY
74SinkPfsTn7+Sbq3mg8SKPWDqlIxZM+6fBmzfsU8wZUjbBLdAEyPwp+eDvUowCkz3YaMT9bGGjy
w9UzoBF/7IdRZ3HoAAi8U2HiMy5T9DnHgioh7WCTbbrNZNK+cXpK2Emk9zptoWsVy2devIFt1+Xg
wUQRVEdcOEuFHKclB+2vE0qXY0rX0R33XLxID/cX//qmqetFg19EVVnZgEmd3dyzibGXIqWkDiOe
YIxeY2ZrPHz5cletIHUigB1Aw/367g73CSvXXU/fwDHj74Ec03Bs1tQvqt9S8F8BIHbYbGXonx4U
ENxuCDUWnsnyCT4wcZ49OEyhIC0ejfEfU0Akz3LTGSGTXe3h8nC9xDFJlfb3LjTrD3KtSuL2W7iW
H3Zwt5WVeS8v4W3exsg0UZg5bUlr0QNceqlJxGlAnjRuPq5gKgkEmuHC3MmqJxyDRlMzN9+qSdjx
w0WF7FuFJCGgMMfIN22H/WMGWK2rijprCeDidgCuOCCERzYodvJgHWbLLiixVydhyZwiwQtFSXhd
FjFCzND8uQh9rGn43z3sF5QJ0L0zTjj87A+PAq9XFcmQDWStgEUMWbQadwjhsj9X5wyjMdL4yI/M
fmw2glgRBOoVCUhouNIZZJ629e63VCEeaord4y3FinAWM9id3k2P0QQrljAHeKNASgmTTcVZ/ryo
rZao7uLYxq8EYSErnwkw4dzkLF4T1WhtL2aJAgQDaqK30lRjPX9IUdvdk4zybDdYPn8D+eUUlSUo
8XvukX3X26wekWQBdpUnJzlrV0FpE1+hAf1NHmsmfYeYW8gQS5EyU3HGAtwrdWvGq8UpGRsD8Hb9
LTly4rMEE6KFTYMYOaiCifvQwdszfQytK+d9dqlkb2S6+FVzb2DCy8hD35rdirftiZeJXZm1rcqG
Ve2DFaEMiG5hRfnjoQUNoL22TZhJQFIvmv6UVHR/ryKhtLNWIj6atw/97BMIs0WqzUX/Wx1cbkWl
DqC7biw6XkVkzGOVOnDtiiEMD7n4OCyV2EEiorKdiqRbpFPfNcNEd0ViO2dbTI3TqzjG6d+xQGzY
LR8gkQfr84PV1JVWmz3BQLPWrg/EVRgy7s//+Q5C/+0bIFWyfhkAk0gkWEsWq/8+LMI4Q9NYMDjn
PrcLiaB8jIjhk5APza/4gIY7J4N8DZzcVnj/0WubD2WEN4XXCP2eZpDd0ndzBL/7R7IMiJUnyCkh
ECNhmT3Zl2SFeeIwmwA2qzL9H3EoSmCfUG1BjF3Ru1D0cfJig+heWSvi29GW2fnOSaEtLXMEX28y
Bjgu4YcebniJSUZAOrD8Cd5qs/a9z9mQUp6Uo7gzZC65QqW5dPai88FY/xiG+5l6iUg++Dbt6mAd
sbEclz0KhAVcr6SHyQfLJwsK2FO6tKeazt3gmr1Mve5avXh5PbtLTivBfkSOyprMqrey8PPhB+Wv
s708iwGgBw0Ow8D7MHqStQusCgnb8N15vpJkM4A4X2RqQxmW7GRDI9ko8U0QoniqLKn4ZAUJt7CJ
VYTQdprSABn/ScjLglQB0CS7qfXOhXhMkXe251zUOZaByb+MZvoCqQagNA9QAXzb26VMSW3qryHl
Bke5h25V7B4Q49k5RCJagw9968YieSZAOFee1MIuOuBe6GRCTahvEzrz/dhKBnrFgCzMGPWPHvEM
b3HxkPIk8x86P30CtubKLkX5D2wEN347xhrxU4BlyYbwZzMcYiqDEP1i6ZJc7xd1G3zrzDlccOhA
LKA9F1ACXkZnTTilleeksgrxqkA7h3DnY6wSYaAAy+3l0ud6mqCE61y/Puw8tDeWic17CbVccQ/h
/9yE9GyVncVulgC/0lBwNrRglF2rH701yyniODhDC1q2Aoy+5G2sFJTdfTSfwseQWCg0LSlpOCax
PPFggBSEmWdsOBjnhY1q60eoiVj2cmt7vBdGmldY+JMsQ5GmZnoSla/H20TGZAtxKrjIukoxs2y1
MwVLXswRr+eU3TFLruc0a77xxNTY4knjISjBCwpbjFh7InmpTMnX1NP9mFxNgY3nQapCE9X6qsF2
avNc1QmDSTqH/8QIIXdq2AKvT0FOnkWL9Q7qAAWF3TFolxKxBC9gn8OMXIp9fsm1VGGXcyxFfARo
rdTIT27isIBsQQeBaafcAEr6DubkORFFgCdCKFavZuSzpLYFDOGoFLAouMWW61t6S7a7W3i7ly3K
JHmSgeEzu0zTuMtJrMi6/c9/KFYfIDeGB4iHiTSoASXRNJYAkrAgyoDGWK5v4H9TXzfx2ehLa9wK
CcmrTapIxn9k2kBLE6V92MlNVBrH0/y1rrMAhs5en909uFa5WQhTaVhKbS1R36BLacHyb/zaGNK5
8wIyjobnJLeJc2ds5ZPC2gg2xSPuehIVmzTi3j7e36fGuUZb7udjefO+eN8IUanuO0MJHPuHgAHg
5ZbiGHWFTGSpTxM0Benz1nM9Z7aPs42iJrpH9jDFlsh7FDHv/BvOJJ23MfG6msFqjrkhW8kQfu2Z
rkmDyk/2PvULapV4XwT6+yy2KPum/yyGPxA/OeeCL9vsKedqaJ5TH4Te1TJmpWtSYjyuXXc9lc5D
HCVTHka9LnMXk+luuHd94hqxO9S1qEKJWqvknhsOxUt49L3Idh7S9JGz9XwbMsS5Av2REpNC1hdM
0Wpjin/CxICtS65+SNovwnB49zwL19M0SItpIzMXZHxf8s6p9EVzXfgpAqMO7VGAfcz7QJx0vHL3
z0w6/fsiyi8TjK/d/Cr8IXSGqD3o1Qyu1NtnSIMD2YgtxJC8224LQ6GA62FQkEGwZGoNCQ94p3NR
qtLACPMY6aY3npgBlywtDlIoUQUWQZkssTpyLoRkW3LetAvO/BLaq6OlSbHffJOPRpYrsXUyhLbX
MYe5j/125UkIEEjAWVK4rneAf3c2N5XMtFcFKzzHRgez8hX8wcRFROpn2gGVVS8+FDfqglu/7/gK
4sGQbH0SjbO+pswrEtyh4usGC7/P2a7i8IVrL+4iTi0/mFFuHU4GtFpCpNxQ+hHfrVbOlNAM/Vyl
L0Eunc1yU5m4MHNiFQRhC7cv/IoGRbgCVlWaVJ5aKSiPTR5j+0wa/Uk1+y0d2KfTCPduf4O36DJJ
z8VFmClE/9EVprMyQATV4pbcPf/5J53d/TG6O4VFrLLSPbEhqTQC/RYDL9QDNhdQ3G6u4yxex/Vw
zZ4eEhedt5UdWZAHokjpE7WGHy4/HU9//O8K5Urb//l1GbDlAKIN3uvRxSwEuKyyj09X2D7fFsH5
laxctn5ei7ihGewTdonH509WhNCMuohSV4FyH63z3Bw1Ua3dHqMdK8dAXzHQkjxMq1X8Jyx1AZwT
ZY5QNim48j/iVsKchcEvjHK1d0KANhKDTvBj8bBUYLpNjfzA510pWfHWrZaxacNAIxsOFSXW0HPg
AA5gGZtBSIJ/NpWGv9aVD6ASXO0OSrWA34RG3DT539bDiOEb5blPTLqOox1ieOx7wgSfe1JT0eEF
3yiVIOBkND3qlvLnpCepRvl7t5aXKUca63xOoJdXLKNbIpB8+yFinIpp4DyLYwRojr7qxmgmRYWP
kCcOsuK3Kf5+qEU6O8GhBGjNW97M4F43w7Hc/Cl7iBFgAg+UKinc75X3JBeFs7bZfTW60m0PIwaE
d1/3BndkU9Cgkbrq6DrFwnA5ZVKtI5GVRSu69Z1BcAMflAtUJw8NbM4vg7dgQhJSkmIz/clGNsal
eiWcI85Z+LhvR32jkIXBaaVXXn8bHhyVoFLmBKwj5y2zXez8Wf+TTy3vKOLmPB11p3DvrWFBE3C2
2GnbZVF2giMvcwOZ67plZWWVSRDcFx+mBCFNupQMtNICWgeReBJgXztsdxhCz4i8rAvg0IKxvsv0
wQN5rPLuthVHObwlOVATv5DFznKIldMMeBvP2QX9gDdKUkjnKuAd2PtKSV97p2bSW5fCsiEptTB1
PUDhQVSm5dSUS/6F/DwqcA9a26RYpQ9j8PItBCX1rPqb7Ps0A9AfyeC2hKmknMD0E/TI7Xc8wUWA
0MvexdkK/cUCwisr+GcoN5v2+sqWFNNBzW2277tjax1oz9At5zgWr08s0OpQQARz+l0X82NHFLg3
vIT+GGLir2CA83QWhQ6SsiPx2pjpAfN/ZGgP6caLmM5r2OoTwHPWwdS+BrEJfx0vikm1t4EoY7U2
8fMywnZFLuTL1DBG8f9t3NqeEG+odrRUQG9iQTktdZ02KyLsauqOwDR0L3tQN40C+GDhK7j/MazN
BtBuJiHj2+TbKM7m7773PV4YEvZBLLXfz2uLbc6b/xT7706Csc1UJvtj+PtXlIeaHXQFriGZUb6d
08u5+X+G8cF2MU4jJAJJ0+SvueYHihLzF9jhj1slAc3tFAysr0F1RwjZCxhUHr6RjCeMVK9gHB3L
U4x8JcVIm5E2ZJuEQtlknTsy94yBLDkkHDQHtrDRb4IKJ8Lo8Vp3q9mIIL9UegTZMDcuXoEbQ8Kn
nJeIvCehpxGbJDElZHxHtrBKSptgGxX9JhDoIcdmcfQdU4obkNRd8/WIaS5XqfGdAdvvXKCkzzaJ
i2YZLJ818PjPvLnNUm7SrcNWt24LRnmG2WmQ8t9u0GdDqbfmLgK31n8+4paNEr937snIzX3hqnac
DU5zw9kj++4JjbIYmTUK20yOvvOshxeQ1SchWYq2wOjmTQA80I0ChkCuuT6oky+ApFoN++SE6XjL
PxRcZCzt/uN9fsAUZUlpV5m4wOr8zWDZ2dTQ4qFWOMXVCsoCkpLjmuN+BIT9UJVrydmB447Wzdsx
8Jvlu4iN7QZb5HKP8/ieTe/wO1W6hXnUZ/SlRvg4Glx8nsFLRlxfnC73QeUAUHUbhw3ePk/xPnhw
w+jb4ebkKxevZZ1PVK4F5b9pX3cnZywm4IeEAJJICYqYJXul4roLDz++KJKdyTiZTH53FIuc3rS8
Nw0a18GKErLea2nmbyRqCmSCqrJ2Yc/YVsvyr0PwEGcVmRc3rs3SRmBDeZjFZeShE3DRvilkswrQ
TayPfADXQmc+bJn7PP6P4X25lfAn6RR4LI3Gm2pbBHOvCFwQxOy5SVf+Te+o5BVu+p6+phpi5uld
HOf2YqcPoQmjtp6LXiHUd7Zc0CpFEsggm+JP++bPzlVZh9/M+dw/DM/Evfz57UITs3n31Cd3bvpI
fVaiEK9Vm9UBSM0OW4w4d+WJowZ3PwktnpWZmUUOowMCVBUYnS7ZvFB+bSYGwJPKfvlWJg8cjKgf
XYz0FKFL5doItA1gRSuQiaslMdMrZdNtMjc8M4DD15ILolb5GiCFZHz3YL1r7SZAX6F2j7d0lDFP
JEdlbXSB2aTntZAcJ1+GADnZqY8FQhsMyLO+K5p93ELqpyZYNuoh2RIxNW9X5lzE41dfI9lYW6RF
z7ZW4S/6YjI6vYFQxgZWjs9an2mTUQLVfGJqkN5N+ONBx86/nvSQb51/WaXGAhy24B0Ta23hyvvD
nvXcYvyMlxwu5hdb6lAs1JIoqDNiWv2BBUC8WnwNdQ1C7vAM88IFc+FprpWic+z8MC4iogpki1YW
NJ+K1OQhET35iZ5O0l8RDq1twQEndFz9sorjT8mGDePyL1eQQztrH9kTWed6jHjXhhU0xw2UFlxC
QP0C9+RyaEByE3DDw5m+pDhpkKsMCGcZ5MsRxqp9u2Co44dMF7K1Px55u3n4EmP9SjLD0JubQyWw
MWgQXA63YASLuhrkU451ofv9jqwPAgW/WG8HMdd+iFQfzdxaTxWapI+/NV/T9/F3ZBLAiaSL8GLz
+wrV6/3mDNJX7D4DBMQLpjIYHRImdldhDZFp4F36PKobpC9z+C/TIgRb2IbWDIIL1UHl21E2yYN7
rbodcVM8e+9vTN8D/YtSa2KKllTd30i4A+v1Su5gMV82RWs0teOUD9ZqUT2nKqol0p5RgigSAi66
lFOTK49w2B0IScgphvik+t4/Jg/Hr5Y1wAkQbKjUfhhHGfwbQxStoYYzviLfbi5n/NLEH8rvA84G
om7a2nr8jC2q4uT6cK72CZiDXywMeIF3X3aBW+QMMZJa8znMohNLQb3NiPLODhBMvRZ1BLd6HPXR
2R1B1AYf7wHEQUlhpM1k0uy87Jp81kpFDmh3JvM/ZXdiBzwUA+gooN8o9M5nhlW6/t+BiTN5Amjx
tPuyl4YNoquRkFGdyFBMxrNOOtW4Kc1L5NkVt/AtZleX7qVJqOjviQzeDeJV84MKYIZSwHHqeozx
D5eIbsYbpytw1W5ndCPuzaclAP+gtkXb5AeIp8olrjP3FY1ba4Ck4GkouYw+x25trb1+gW6QrBej
BPcsS+xjO7zOfZRtWMvTQLmTUYlKHd1Xkc0lPsi85RLVfZW1jkNwaBBITfW0KHNwUt9Loi7Xsam3
UZ0vmmvtVYyTOZrhRHiMQeZekhy8d2nrVzhQmRC8abMTVEiIvCfhqXUG4r1RPAY9E3kYjcNv84N8
4742FWlqSMBEJzlEPh92ClD7hhY4nvf3+hKFQbJLw8co+Hlx20kuSKD6AbgA/apm4ENwavfz4tAj
HbL8Jjhii/Rz/IIW+leZu4gcCBwohL1cSMgaFvODbsAumLG75tAP4dFp8DRzgvsZC6LBowQUuLuP
w5c15wJ6GiJo4K15QH3W5QF8cm9b2YMrK7G8TJwmm+Cap1JYaYvLf6/2Xw0vk+9u1iDAb0rV18MH
ydf1qxczy4hOWnf4e0lf3Ro8CrGwHsBb53R54IK/4XTUoBy1rM4dhU0EKZTB8lpUjqrZjIqXCXb/
RhRuaLsEsFJL0+79MBPtNya3EH2XGaNgGil1tgJXVCkoV4inYTHcG6WJKFk1OsugMomT105mnkWS
yPpiYSobW9Dj4E+TCAhfhAQYVqXOrAqdGU/G8dSp1MKRmANHHZKxOSw8xJNBMVNNw9fz7vyGMyEK
oEOqceVkY5m4EeMX8AaiAS7uGB48h+NvoGGDAC06ue6HvQGRq5mjIpZXZdE8aI2Um3F7hUbymw3c
bLPPONcoUfku4K6gUGkXmFeYmUNtLDoQesegOZvvyjdLv7seQpUDondrIxsevsUfxXzCn2Tttg+t
shNpLvX0uyJB31ZQT9HTZ1e3RBDPx91+wqkK7gsOoBDCx8BOUVJMR2C7E8bYT/TZeXdawJ02C1h4
qPRUxGKs84zvRpU0DEHtLnYJhJfDiD8Wx47pbkiUAxfNMt1offrp3POFubbT0Z0n6S5mgZCgRl7n
HSIabOFG5ZcXxCZcBqQOKUePdMn4RqAexyBeoIvw/qXgWT4bHV+cign82ZSt/UzxLwenFCqYi77K
hSBfA5UxPu3dibmMbFJI5odP28wGPSNhE+bnW6mScccWu8b13DKCrpx74MbyQ5317qkSSvO+435R
zoklZXbjQmWw9GB2Dvz/KQzgmz7qP4qoVmmQGqbU7p7LgSO8M96sarEbwDONjSMGtgra8zYJrBV8
ltukiHr/1V6hhq9WZJ5DtqfByBq3rUfkjp3yfOFAVuPrNzZ+NKvOVohgz9SOm2ubUBb27iKJcW2k
KbCrSfOg8KlriLQhLke9tVGb6cTqjmI0dlZh+v+2waALt0QelXX5oVrbOGn4AYORGAOSq5/DWywt
7fVz05Z63Vf3WZGS4Mv03JOaedS1JAVHqRXrz/TwkidRvk0u8UOX4lAwQLitHp4IbWA4wCUEErpG
Gva31xFR6g2YWaHmd08kqVP7c7NnLEBr/dVFn1KoEhRK/jIgKYoXgX7JfcpsblBSHSa61xetfL3+
Q3s4FEMsY0MO5cz/iGFdJzto/5RvDpUzbvZyWDQ/oi/F6/yvq8XrN83VAM9qC5uzl9K6r5TOW4f9
kn1tiSMHio2j+h69OLfYGPigY1rMm5ypKzObKSQLJX3MIQYIRdGSmSD4ilw5eBRmS3TxJI5JbW9w
IoTC5bYwopbfTxZ8Gd6shhBgxvfKEHO65b81W7mCuD9C/BjUGyvlb2pOwQ8tmt2O3W2tFlR5GwRh
nNlSD7cZXQNcvQt+xpSVHyM+6Th/ozl1RpIH8QmTq5CQ6qWefbtQfMn+1fihi34rkHkA250lfWG8
sCGyOELkNZQ8Yqk3xG2lmka7irT7zjox9Cw0jCpEJIMDSPSNQ9ozQgw9Td1zAAqEAVFvpnx5ui5L
PPM6wnwctUpLCesIC6CU7OnmIfrkdUt1BaYm5+NsB8rWW5AP2XSK/bn+heyDSLzzPE6D0A6U0PY1
KQgOM2QE2fLS4M3w2XqhGjHv0yJ4NndMvS8IZWCowJT1TPNgy5RtP3OjPu30yqJdaHr6CA7SMbtZ
Kn6orf1bATM+WW2SJW72Km30T2THu9ITzNA/7EyQS3hLh9bXYgT9RC10qTM3+sKN5SSjpc5qW3P9
tDxHlQx2Qd/ZzU4nYKukrTomwMBBy/KDa9B3y3mGcuRC9di6Tx6VUuLwoMj5uUnQ5dYFGmbn2O2t
o+GMTg+0tmFHVEF5/iB8f8re69E83PXM8hEN4cexoT0kGVXp1PbUyjHS3IBApR+TvTnaL985FhEa
dIdAH3czPlMLvSWMU9iw3dmexFcf9rW4LJFKfR1C5JY4VQSv0auPm0jJ1NeWU2LtYC18n3GkBU0x
MFMBhzAvlKFwYAUisTBY8NsUCpggfjbQddIPah6fPqcGc+iwasdU2iTtXgbieM/YrjGtZjExCJgm
trOkMN7U8w/fDL5lg02qADGLkfpce+2MSaMhxg0/8PMMuEtAPA4vBhCXj6TGGxwCVYYy5GJEczpo
Uyb9t4USIY95AUm6aj1rn+Znn49jKGBBP49OzKjjznFje9OkhQqMa5KgWZZoKwJi3+Tz3FTO+2d5
H8tEQUFiVKnZsbZtTEL8YZSKacYdScKttimGGgTAEjAgUaGtfJXJWYepuHfchvZqW8ZBvcWnro79
kVYbfw70rsrXpRlrx9NvFqmXd+7mulCimM1nA2tjV3+1SdCvjY1YEf32nepkmqkYRdJr3rF5ds1o
x39KDm4Xk8D6X1kWngOdidJ7oNSn5RGJC2xS61GuUvURFFtM4PPc097l09nom3Zi/FyzvAfznYhb
7GqL2JqAUxPRHvL73I27/dQAJBLEMWNYft6yROC9Qfay1uvpNYqEZxkhHjbe0VdzYPEWfGRZRtPi
QPcFKheWv9smimiXVATQsgjjnMUFQ5CBBkcSIabENcFFzjpHptPEUIB6ouV5fOpXJzF3HepvtbAk
/BAnv2R71RfQMbKnzD2Y5zR2j3PTrPnyMlS1JqQnH925Q4GHVU7hL6An5VCn+rnOmx/FUTivYbQP
zF1pzFTCVY5egfFLWSPyxJX05jqmZlE5vCtiED+WVylhH7VaR66BmHssKfOcgFhvog8DnEH93mU4
3BafsV+U4tZEuiAkDyyVpJkrzuxLOp7Xgbg6fnzrBHgsa/ljTkmwNLrprN50EiCRnDuC8/33dq1i
/a1WbQ4NB1lJGvkjOtVNXOu2u7Ego/ppdTt4kYEKYHt2fokPdvQ5Rn6sn0n1VvL3zX6z4PEomKfy
/KzpIxG/0Fq4L+fjRMEltT76BCq69SWLq6O8v5pMxue+X1OnqSlZigFn+AiI+HDGy/spY3tMelve
e2FfADxidCGRZeQm/537RvghZMS3iNBR15i6VgUuvwXefSt22aknopTSBshCLVLCtUHogZuELCZe
jjWG093FeaWKQUQvxIdNQSwALJrjYf+2rLQykxBxPccz+IeEBTpdj0JYBtx9mdKjJCI/fl+jrcBD
k7Vf1aTC+tMqPMXPl38x00BbTpwdbtrGk9Xpv1zX0c3KWlVqLTcLMBivvmmpUPteF5tb2WYsBzP8
dYxOgE42xLefQQE7iiqNsKcr/9hBXnukc/zMR86UyDjoAtkgkfuoQQxlWZWDH6cz3yITn5ewAWIF
MhqWN1wDs0Myp1WYEqwtj5+AvTwamat7m63Qd+Stk2BRZCRpWuPAoDe6O6k+2p7YRf1wvNe9Rj7y
9z/G7/2JBI8EKpUD0r8VpFcBZmpcBp5YYfuw7E5R7hHRHQ7hWuQG4E61wCxVAasd+shGK+nE6/21
Yhq2b+kOf8XNf+dRssgwSXmvfopphw3pAENn5xJsDLNWDsBZdaRsWC9guF4rVoqaLKRdBZBGfr9+
DDO4Sq/P3gtXfhwPAB8cA8VMXGR+5eHmyfNzjS3iOP3bw1vOoOb1Ex5WjBZ+D+4rU6Ov+MChEwug
7ozFaSvEiPe6z+dXZo00WEMmjaw0MTPNBgrAP5MTfAu51yL2BiUwO+F4nutfuH+A/fdcTNQMI5NI
oksLGxUm2d81jo6VTtX21YWfSlT++MJuqBFMgB3xc7Z7P2lpeHkclQt8q4yp4Hw0BmVNgA7O04qw
rNGWl5iH+YtL1vWlyhmmCPrw30W4WD/9rRcO3lyy3hl6mpygtkq4fVISprsqvRRVphawy23uGI+L
taJMQqJTNAHnuNeFdrtBkaKjq62qyymdHmBeYEFYwZ/kk9O6N2fAOmutnQ53Xvzs7VcYO9tCpp9Y
5XYUR2MYNk9z9tGGbcBqYt4a8V9rRWQysV/RaR95Ll+dVze3sK9pogfCqoqPD2qtSDY8pih8uJSl
hC7BcMHNlPjUx7W5NoqSwTi8i10guEuxA/NclWqbKBkqhJ/sGhvqWmuNpQRQaXimZQCIurHnk53h
pJbwyXC8tCXPX1z6wFQZ6agi+boeZu4lJ78TLxz3IlWaBbVb7mWoA6yL6X9bcu1a5QbnSsVqTjUp
tbnTjkwYHJ5KzCMd99WBHd2DDBITL56t6dmdbuktPUoIJgj0FvytNcYzXCWIGRgdsC3+TZQ7q6WG
m4kqlwcwpbYJCDzQO8VuxcwPQ96YcrfcBBh5TKJ2glh3G1TsJyYG7c9r7y5BREbNjqBob1JbtVI6
g5UUsNMBlSVEDc2cxWisoRVcC5UZqG5LDd6ds0uCT/SRJaXZPjLt+U0C1T8c/FUGTPEkgk8KTjYJ
FgrXAdrSfISrltIeaqVlTCREwzlOLaK+rzhv6APzB1D/uCEQ+joSH2ZGieKGU1WozVzvwLWz3DH3
BbOD9hctLNeHAWqnLySfkE4KUpwjFUHHhknUxkrH45b38XTj6GW4Wktbj84JAfMooTk7iE58lUVo
EwYflPsG62gO7fScixBwKOInyQuwbW/KmKrjCeiUazE92olvUwNsCQ5nWoBRGtMSNBCcfBWABMm2
JjT3KyNB5+Oilp0w/Wqv2nC0vVftTpcih9yUrvKWQOuAZikhBxYDTlvzht0J61YTyNFj1ngRgilI
o4tegPcAg1mAEhYw/rQrgMVv0El3kYQxKZDhrByySO/l3lNlb9ua4LRN1PufKb2uLQkkJgGhu8pC
iohHg1gSPsj3AoyRGyg/Unit8R839kU7evi4LL1skeBQcVpl2Diei4QN10wLRTMaKhMkjzjrJ68S
zXWQpc4Keey58T04zn2w95j4FZM/lBNxEhi4E7qN+t3QiqI0QKUYp0mYo25KQ/51maqKL0w8mTYd
1VgSDHQTl5e0DBHMoLHKwXGuWNfEJvO/OJg1qQkkOz9HJHhNxBw6zBqGDuUFMpwP9QRw2nY0nzLm
WTfpp+Uf0vd9q/GCk1pRH37LZlLkukBXlJzGCAC1VYegllpdMyAefrQCISDpiuqyxJ4dyVoFyVVe
kYbcdeqTR8OzmspDxR32wLyQbIBsCVXFGAFVngEajFUj8BC/4ww9f/tQQKCwaoCKKEhPxdV31m3w
lwtApwTJtXs/G62kpb7caqpo5c98M3ePu/47H+lv+7/nKXuIEp5pWhx4prTHO8rlt1f4Y7fXsJNv
beXjHV/an2G+8aD+aQ2UCdW8n9LAyHTb7bI2JSKeD4KpADtAIzv7/Ojwga/Myjw7a/ILHx27B/2U
ei1txURP2LKPiYYIznrzXVjFSH0nmDoHymidDM+cMt/zIspdg3bOQT6YbUhic3FLmIiKoAq1lQyk
inHDIwFd/GuNTDJdmGH5bYfn9nnEATCTNFI29RwU8ZAPx8KTQvQxvQQN1wpgonqrM0RGXcEsTYDI
KNzfosLoP211fzpRtpBkZeS356hDaMq9ArWqILlNo9vfpgdnPTLikH6MbKbZryqO0RMy8tyyVwuX
zESrRnWWo8qS4zsj3nwxYdOaG2uQJHRjPpAchzKOKzxHbGT8UnXs3h6JMHoHbHzWPtifdx9fRrqO
VZBIpy0lgDGd9W6Ao1c4c744am+SoX23JybO6kMvXur02FifkniWQ6inopqQkwmcFVCLAEAH5j+Z
Y7GRAoUVjpjkNhcQiouaUtGY0Y8oe6Qw20Nuvrh1P8+ziUBPf9hPqkfSjNWZ1xB9dAA872ZgguPq
ZPthLWEMq1MFmutEpu/ekrHUfFLXQoZuhjbNZAFsiaR3JPdiLcpUnOUsBmDQHCxUUTQulE9Z57OA
iDFwtNlbPZa3OpNjZL1FhXRs3gKgfBUvoaCyOPQ/78+2VhY1yUt+uKcHm27gAP5Yd8uEdCYOu0PM
WHA3hCiU/8X3GWU5/UmtplDomDpzZqdG4dscpiSvCvaSzaGGvbdOF+R44QxlRT1/zDm+HBC/M9hW
pP/LIS2syd0c0wL87bL1nci9N60L6CUlJ7sBkbNAI62X5/2fU2N7q/++9+maeQx/WOq2zFR461Pb
FnajetobziLHk0//AltXGVTZv6yNFYxAA7xm2vnbethMFyrI8fGtgf3FY/2pzlL39H3CbQ823uo1
YXCjefDV8udTXZw7ai7yMUGKeZrMvxiKxm6f9ZWlYFCZYiTMBeH8H87Xd9Fn5xlfTzRnRafGWSS2
hyNRPEbnUlii2cyT09u0Ub7ISDEBgZ5SmSl5DR4CWEfXVwf4oR7YBQZQF2QOPqvQiPKEyojA9iwf
an16S2DVnOu7wFqNvhNrAu4iEpcsCMTrxGXoMwENkHnL1BmqqDDZ8GikyAymQsa5pj6Devj+f+SC
XFJ0Dj+GG+u8f19Z7scNoGqPKodhjQQfZJF6B9BHYL632OXaiUMXs11ZeRB09dRkW2rfabNXzTjH
6egUImSZSTppqndJX6aT4cKdufCvlznu8VvFz/spMrETAEzZSgkqhG8PX7yfvcmhzQ/HNXKqtAkq
h4Hsg4hvFb7eQvHR61FX0E1aXBicQgKbPDaDVb13mgylyQTJKh6J6CA96JJ+JJapNVxAd5UZi1i2
CnufiqAzbFhM/2pbbYD/HFNpC+mjSCy1ni9aL7R33GUyP2wrMO2pJ0Eds+ZUgqNfGY9NJ9l+9ahr
lAF+tPBxSX1TDZ/+pk9iyeyS2t8C/fv68OMvEV6zyAVbghvULG+5PdgvpKMxw02LPJNJbfMibTbM
/KZRXUH0tsamEYRCsSzHeAf94SoMPrlbbRWdw10ZiD225iJHbDTERucLV0Iuc34+6XPUxI3NIBJf
4FVNTDxUbCBQqfwXyvv/ZIxU8bpmX4NnEEVvLE11MoZy6nGh1gSZoBzRxV/42LBLEE+/Eg/hsGj4
JC27fFuaoDW95l+36LgEicb5dc5uCKjrKp8r9jH9/RiGXL4ROzaMJzFHTEN+l05Z09wjnp/BhFWO
eWiC1gA3vK6dZ9SaJnLrj9d+msztgB5VSNA932Z7DEP2/rk5P2C2EhVPKSlnHniNSwbTI5PueYRu
x9DnXp0rRCYAcyIb6ZuQEST+W1xwZ0rftOWULsq1wIsvjhXnNGN6XPCl84CmEsjjyycz+Xa/00IA
tD4ZuamqidxRw+5of9pAx1JLA4a8roeQoo+cB8gYFtSGSPjGumbeQ4UJS/Ks5UDLChr7GNpRHJYX
y4d4ktBxoXdzbkrf+y8b835KEs+W7hQJbKAQ5npQs2u6vHGEq7k43qMS30TFdOhBS1FUi8rUh5z0
4s5T3rnrDkDMXmcYyWJEG+0iWMjPYAJAqCvDK2OcnCjiCsp3xZ9sqnyeRh/wp4A+l0kTgD9Tb6XC
TngpaFJovXYNHTtoyVU9rfxirgAU4a/wkn3oJ1tvg6/uX/NPuMs1Ku/uPij2gyliacOJcqgs9+vy
bfuGvj4U/Z465DglS35O1fhvmqtIblC5QmtRpy8L62V0cLtUr11bw7xLvylZUCO8x8NBsPrrWDC/
EgEOlWmER0pC93K7BFCIpoSAJv7ZBXbCuMqxcLYURtvFww+TilmnWojjfWNPsyWONOtcIFx0MXcn
jdOA4vaaGbS0zIzEkNLWJQKrM2MrNTPMvVn8JbxvN1dZzsfKtqet65mGz/Zh4BPp8MYrKxoZAkDn
/BYrZWkHscV1SlZCE3BjgFklPwcuaorRgWPBRS3ffT6475LIevaO6QFa51KIhxDstCbkz6fV5938
xBEGaTjwENl4jCkglekUkabCFnEyXH6ZuKvZ0zY6Y5BDVAqPUKHL7xH0czqNqXz8yvnmOotk+wuI
OwzJef1UcwAe+FtHkkduAPnIsc7UZ1zDfniu14NoarkiUIFRam2iASEw46+XAXnQW9v0ylaExU2B
f2vsoLw0/E7gnG2GZ/FTpiTcg19lj/JLljq7SksiaY4qhJCtpKWve2zzbZMasmmayg78SP3gKMF6
AvPjkwKVqV0QTpQuZ4aLkB5v06UQN4NleXZNcMaPO3roCEZXIyncQmX3bMuA+vkkeHgT92ka/sQX
1AYJ5kRxv0pSPsXMECgCPGwUMYF5/+Nyz+2InJ+UMtxbOX4nBCb4I25rqqIaXOm5Ya02aq95Nmzk
9mVL6syeBvJDKO3iiddf7fwIuEoIM0yxYyY+RUPvzHNBqo4yMTiX/HXEYURBOIC36p7BzWiuHo6u
5Fm4+JATXK700lSyHrlWFqFVTMCbuipcEJ73+vK8XVneJzW16wp0gWSoAct38jfzQElTQGKN2DsS
FfXZWKlulE7Sl1WmsVXhuPYBd0TEixtMZ+4KtKQ2mvPNrfUvyicOEuDXrcEl8n3JWCLKN1leuvyM
wzVy2QH4WpJiAOerwldQHltLbdWYz8AlaYFmXlfCq7RWjE6z7jyHZeffuuvYnx09UigAlJiO7CIj
h4kzXEdW/jSbHcrdGLTucjFLz68vTbRfV/pq1a7gJk+q478XteNT4GYgDNgCnKZoAg6a69Z5iS6Z
5ENXJfi+wzOd4RR5gM63wGPBu3VvZHYMvSCoqCO8p0aDJla0piK6UuaQdII2XEvZMmJQCrzokVeJ
sS+8TzwyFjc8yKp4simI3kqRtew1WINrazO4lX3JP4Zo2gXomVbGCfgfKh+OdJWr0E/iwBtSUoo9
XZRZ4qHMGfLOlUBRpycpOOLDZKLm+AJ35fnk0rcUQA0J+8odpZ22sG+awUVc+KQI2RmpdeoN4xdQ
fGj2mLrDKtTVYp6W8vPEytny4eNka6jUtv1fLnrEQO/jwVAxGz2VgPTRzmMQ+r5s9/T2iFJu/r9s
pm3kYSjqe8vBtZ6tLl63mCUvk7EYkv49QSkHav16VkQUhUy6h5tk6CnXKAn02Beo7GARjmTIjZqZ
SYi9Z0On4yTgjs7zoP3mW2maP7GOQx/SqG30ggcB7UtOCfxfINyXf25P19O/QIDiDr72P90fHUdq
BwhKWLzan9tCYpmqcP3N99QHEbXk7pc8TVhRdmJJXDIr7Oa3eydI13SgvcmIp4ltPm9w78KhH1cV
FaSmvW3IoRZnmeUxdtYW1ENbH+gG8w7pgTBI3o+Jm3MtEx18YCWmeUl+delUODpPcgPoE/fI0IfV
atcPyNujqUoUYC+aRiqlmY6MNwexTqJHcrNqKW6F+FHhzxgyehlhagL4rm92An0COFeF8aXMLmsa
gN93wp2ZNbu00/1iaYYAt3Cl8m9Gx7D6KfKNdbhA0e2SsS6RmO3ytG9wbNtMiYAc5UxnDSSd3FYN
wuzzWiHg5EnS+Vxx6WxFC7qCCN2xTaKH4gsQeqY83bP93QQpEYaaep5TtA3pFz3KF/FrW24T4emX
hfH8E2hRlDv5w1dO3tAYBewb5yt9GJ6Vb2QpD4oYIK7Ys4PBihby7KE5yUeagzyWwfnrTr6Mdabh
oQ+hnwiGmYxFBGJrHz3d+VUeVklaJ0Adhvo390JUyHHhmZLkwBzNRZSS4VFH+ebwwnnJjIArdlTZ
YASisezr5g0FpzPbg33lLs22uLmAfIT4OlfhbAQVaUwYjMiqzXg2PDjgjalW1TFmNs5RhpG0HsR2
wAXmKZzgbTMbIL6ipVFPYewWkj1p3dsbfwumID2wC5w/mlYyLM4ynpce09jR7J93zdiCPrlSJzlk
8lpf0AIpsJ3VbKYLy7UAFyw9cf+yCQ89n6XPOEQsu/f/4w3TLiEjnqPYeN6A0le5TWR9l/9UCz6F
5GzzR+KjVPsNrb12NISBgoYnwGlls03uo7uQdyu2hllg1MN7NhyDOSvC7dq+SOX2M1O+mk7n1Eu9
raFy6GWotkauFtLQgsRnOG6nR42tfn5+Qj1AP/l2G3oavCOq53UpjfPk3waPM3Ey/mG8zQtmYbe6
YceWw/SKUd2nyYssOPPFZDmqyYgJFzz794ehXCnmy18Aj+gbuzXInUsbUqiXKMNKt45+zzx+Rqtu
ThQYdcuMGL3SIvaxU9k3zQR7/UsGJ7s5S+PK5j4O3oZisPrMmigU6UVy6hfzJtzOAh3VH2RgdpQn
S6v40H+l60kjWbbqJatsiorXuyPcYffkQa3H3/GpR+jg1/j87ciHWkffFfT/oQV4ZAiAqB3QYaQd
tNd8caWahBv7qDIyd3JoD09yqU/JzuZNxCoa1/Hts5YsqdXpLeJbsabhJ/shNNQr8nNRfk8miQAA
Pd29DH2YolpuD76kcTpLUuEXoGH1ONbpLS8udXveuGyD2VS/mc/QfObiEVXGOsYDrC5x/snmY1PQ
qtroAfDzuVlkrix9l4vsr87s8kn9IX6mVoiTnqOUKWMJtHc6d5ozTJXFpXdoWpltRLthurGAfGUh
JSCzUyS/9sziGBAYa4+Lv6UlxgO+9mwKl/pAek+zFQ5uDCoaw/qBy88HCcj0T6RBRgXXF1DsObDl
aF01CvQRvvswhwXHeP9Zn/AAxNxbP2PSduIpzXG0O75UBqYfQvghfa9mmr0uj1TI4SRc7MegQXno
0rADJdQFlq27crdbJHt6EXW6l+nF2z4udKRohyg4k8182GNwbCHL6EgdtxfKfGQKikpNZ0jStRos
GfaFBXh3QNEarrRArM/2H7EVFIoRRRLqSZI3ultXuyiflatY/ItKEB2SjU3YWdN3yk31BYfH5Kbj
c+4Dktz+2ZvQoSmTASJoi4vvJFWySLw1D1NjUN6BHgVC56COBbjWfWfec7AtwfEo+UVm+ZSl6DZ/
TKPscbE8LtoUVe/fybf2l65mYf+XwB0FYN3/rOns8tKS+g5/ErMA1Sd3qhiDZspsz98uvHhi1AnV
pf5o63jQpfKqxMuNr2mFN6ub/4/ZApRyTZb4S6ETxpyiYWhSgTBqSkfSiCX5xD5G/ZEL2blSu4wC
nF+dOZ8MKWWQyK9CYvNrQp4DCGBPPoD/8qJDanXdUcw3lChZHqB0gnXuEipFtHMzyo8iSldkWYwN
Srk4FRZP2JCilsZigIgrguqu9RJ9m7vrV89cU6Xz5m6F5a2amomb1GlZNb0+zDGvnCZrZclbtiK0
ik/Ge5bNN5dHKrMSZPHJ1FoOL2EujM0eQ0ewlvsnvB1772ikj3N2jhVeW1t5Gu+sWjpIqOR5/9Uk
+HeRdQQkyvOL426sAuwEias2n1g4wAtFQKuuD4nDMx9tme2fi3PbG6QNTuHdwn/NNdc90zJR2W2W
9rpDSFIg/cSySmkMD3kNW/tPDsT5XKl1WfFo4krT8yB/AdySCdnED2uXrpZ9KYgF6mrR06At5f+8
BmEbENIDUemHCSF7+WcuDzHwldZajyB9pdLrIDpE+e1LrCSN1jGpuB/qsZZdB1dZcovkEUR7Ii7F
noVxsF+w8Oz0voUk7svAqX08DIh8OKPMJ94Pe74yPyf1DAhMiP5XAtmd6RXry2hDRsPyQxmrWoes
T5g/3Bi6qo63ghynRs46YC7gg34Ah1REzovTbdPzmUqspZnxtgfmmvaZ9kda7xx/vVPutFoxEnsU
DIJhZVr9NmuIz7RyYvxuGUG/ogSHeJnfI6EXSfcdIl6V1wm7OcwU4jievVj6EpZcr0cr7HYitkBl
j5Yhf86TNCia/6HYOfoqih2crLbaWRrjHxwqynpAJiSvRUpDWQ6nP9B6GLj2ftRVs1NLuvJ7PGCZ
h3GtOJtzz/kSfscQb1JoUifBlmxbwZc0b3XufoDL625zXdQGDlNXGzoHKqN81YD2W2WdEmGUORGy
nBBWiKqi/fP7vr/FzhbxRR/GlZMyGrd0QaKPNEoKFfNvlf5Klml/x0i4oy8ASW9hnfNjZcIguBH4
YX2MruVPvVYbSEAVC2nt4y3R9K0pH+EZHqxYDYTf24ZEXh7ltv9j0hFlC3hAQx7nSD1AOjeTiVxq
DPQ+Qp/DDLD4WDL/5AsK2B4/Ybbr33zkpDMZC1TCDAwAfBXrjn6vvQ3EwS+d4ey40fZcWBJEq+aA
Hxs3vSyE/IinSEpyvE8wYONygAylSzwugTile4QNbCeU5m39Km6c3EtISyxUUjhsOzTDOAvwtKZm
vpolX7+oKm3BdlNdhqpQ70H1NpFB1rO5lMdhOgGiQ/RhvP/bHPt01hrLu44NbqCLkdo8SHb4Aw6M
8w5jocp+B8emn+Fkvv6Jl5xU793BzMBmmLBRxOzmk66/Yk3PSa4ScYKQgm59JQvPKDl3X6bGaEtt
YP9LEDv2JDs4BW7KGTPlq5aDdUbk3v4E69EORM7o45gqn+4lBNpflPHLMLOGIKwOKSjo0PCY6owv
Zkuv2m9pu9KWk8+/XJZNz4bdl4rjfKG98t3pzsfpakBKC8FsrMCgDEggLa9ZxYRyUipJ0la2nV+4
m5uKhsIZohgSrGb4UG/XYBRK3z3WLoa8UeyyeWP4QqyYSadSOQxBLQPtL0NHlDOci7IMwL2l2BpX
NnsvVcSkEuEoz7moRlWQFua4u7GNBzSAba4+SredRibT4km7H0FY3oCNKpOjlkbbllMdlPBSW9gU
Ld0Y3iYGIwCg6qD7Ei2yYtf9MDmWf0fNKZO9q5Cq0p68xNqyx6FiQ8tHs7oDxdjB/yizp3Q/Rqeo
ghAKkvA11SL8NVuGK9zWl8qpmhwNb9A8xIWg3zFa1ZO1evACnEKgpsUvdF7GCwsUgWmlP41yAwyX
nDe7a0JZItfZfIQm2SEN1TNvp4Zd2YpluAYcSXDutgQwuCfin8lmg5LK99L6dl2KkRlUirhJL8e3
JTWMZfU+7/LTl/hrSqOLTg2sH3t1beQ2kHHTX/2XoZ0RmLMoNVkrKHKGCiOxu6QWUukpBE0dcHfW
3M+sGj15JEiKzlJoQ5L8cvTbubhfAcDvA8YC23ACha/8imtz/6tny+BlI2Szs7LJNVQ3c144JY3E
JC4iWU4zhTN/5gd0N8cNe9MLyOdYaJeBN/VkknwHSU/Oo2RTUZpIK0QKYckPYpawkNu0JxLdVM+1
nOSY0yLGC38lAU2qnkCVlro5t3pKpnD+IKXXrbTv6iE5arVH7ZWlDboBNK/rFhzEiIuLOfdb/wx3
N7nnj7H3KRXOFy8IgTwrFbgTOZew3eyRoR00nYto9yq4om2MhH2/XqelBPkR2SStbI9vYs4WZIDA
NgFFXml88EKMx4lhNDxdj+LE9QJpmxUnb/gj0fHZoV1rlg3z0fgX/ryl9rt8dpsCFhcXzqzQPylU
Q8wxtV4eoAnSqByX2VX1s9qiu7ItsBJW5aUsBYQMEaR7f8YeTFf2bRpY3x0ZrtAJoG+ON/slrAHa
JEyMKo8fRoJfYA8CwTzmMg1BkQmhD4BT1z4qOzgswe4CD4AKbTLICbTTeox0JxoWWNElrKfQDOhu
ikJrfl7uyxs6IdGwE+O30pELw2MyNjrD2Vl2Qmih3GSzg9sRR7xs8ieKf+/TDZrc91zZMRfb5s+Z
MWsRQksyEDpoMRE147vfjG/+mJ3dxdJ+cFMv9eM7Zr4hqfwzOBrOPA10XuPVpre5ALSns9JVZztS
uYjAOhFk3+A4TOSYF/Xpqvk9TzX59GUvlZ+6Yxiv8HecXpXWxL6BKc5bZgFDW/TOVng8W+K7HGXk
fX7H0Hp9CNJ/MCfPIHjky+kaVfCQL8p1hbYVqkU5YObNLlrTwFo3WG05DOw3Kt+1VQ4QMHZ56IcG
16Jsc83n+tL1jj/bW1P3Dzzl6YaKx42qNTQRcMcUwt0vTcbeeL3jhv/Y5Ko/v3CpWKebE3ce91cl
PyMAO+vzvB6yA7cxLLm+PeBngL7hg+D9VIp1lPUZEE7kuOgKt7V1pX8RgtR6AngZ1TDg/uaVBMo6
8e8TNv9k4GeXSVlF//jMfziQzdVbXYNnPLzgnwAsXc3LjNCuGYm/s39iq675vBEeCn0HvbX3TO1g
niEcl1PV5+FQDmD0ewp20EZn6ojBRGzeusb14IrMF8gniXbIeTz9b6UI/0Z2KuB6ObMirweu/1aq
1uZ4RFHB2H4TXkDBHRPkoKLEZNxRzKH5TG2JR1bVlSliYWiQe4t8V2bkgIQeb9Ejw0rkPKJ7MWfl
rtB3Uof8VHEVkLa711+kMvuf1FIlGs2doLB1l2jvm2ZqHBaf7dIQZKpcGkuTOmz/Ito8zjEU3cG7
gZqas2NJj2krAOtn999atTFp7NAHq7CJiGwBHFghqlKWu0/leRBIY5PtNcecyaf8ccnZNl7Gs/g4
vaYjx6G+9Xn0ztx6/ZDPpfDsb8cFBX+UJhg88CFBBNPTDjmdDptiUyFhraiG3rAlu4raToqqGIZs
XN+JEXbNGphKtRZpVqnIAz2TvrZrlvN6oQrNglWw0Gkm+jcBkDeSMnT5pjhqtStu7v+TP5N1pt1u
qIXcGEe/XZyK/8Bb9rzIHObjxJCB5gHqsaP/yrgBSCci/v/C72iF8bsHeGsstLMFL22/JLzuovJF
9SfS//jpywDtsXXf/I0CyCkmjkRCtvHp/Ru3rWaS2orzyaCno8s0eR0+dbLWcvASDsCo6YLVsdEH
GJbpMpQt/wiceBANyJPqrs+OYVddWuZ2LPAXB7LzCm83ixbsXNKGxnH0vAN89h7NqbGxRUQ1ToaG
0bsxwgvKEuQawMVZRvBaRxh9f0MU7N2Bt6zDoGG9YBQ58Y/TqsYzuqU+Hd3/hpRRXkHpJryJPVN/
mjwQsrXxmnwApmtC+HqdogERb8A6B4EnFE+ABTgfxXGCO/DsccHeNwjmkK4xzGUvYur98VY5RFsN
ZKXsZW0xooVHjug6hNdfgs0DLNk0lZnYwoO9rZNicand6n2mWvts8q2BwiQY9B+TTYPFLR0OyFcr
05olll1R5P2VacCgLatmv3Ajujbq9v61jEWhj9EHBFS4bkvSQUspjB6H0ZKyWs99JF6ktqWzWNJq
g2DOCqtJ8l1XW30Q7xZ9/QehsCGjoCDju9Zim0dCu914I3Ndzu11elQTVf2oZgtizuB9fMxHav/A
G7fJvf3q+tsV3c4BstETW1gXCNit0f79RBRJ/85p0dP9ElJTlXoJo5WruZZAb4x0nIN/TN21fIe0
JfoK2aX6R13wJAglQ/wMolktJqbDr33p1xdF5fW2OF0VaLakLio6t1UkfeognvZId1nbeSuJgRR/
3rxjIl32vmWWpi+AuS/JL+D/VJt1zEd0sd1hfNksQ3LiiSMI5Uq+F4g1WyS3zA7SRLoaTfztorxt
MXRoA11omzTXRkvS84SWzBPIi8sFb5e+EP3hrZ/07rdAD7fRzrA8ZcIglGrd0slWQeKkG2T+M8CD
dQYoniakWFijYNst3baTbpwMmVQ+ZjgSI1Weh5b77gcy5WbZWpsjm04xQeH3m/hb7eqo/4AW7/Wv
r13zEV1bMKKrHsQqkvWxuwuo6IdYWc1RSRSRSAal6fO5VUtktr5oup23KTQRDpQuJ8l/rw7GIMHX
U53N6ukd42wrBKZkTNZO5/t+yQbsvRzx76HwDi+Sr4zkIFNr3PHKLKRo8Gut3hnp/YXJzn70vHD/
Z7eR69PLEa9ZFLywcdHaqBBg45Q5hgjO5bk2VAaUxBs51B0Aa+WhI6MV245s/BCpWbgHyCuLCYQH
45VSBB0N5z5IRrhs88ZIGezV20XhLank9FLpXc6218pkkTFSC5CcnUlPvAuQpa+NRwDCCLA/hME3
3Pre9Iti/fykMUWIAsg6z+72BOiZF9HzgVeTZs4lBBIula2//Gq9+8KcxJiBzSF57tjEKPZfinjE
m12av5w1CcEuz0J+9nGMEa/jRlcW1to/XwJQiFdY0UuOoN7r7LR8cjpGYvqT+S2LchjH8nSlj/bC
mWYp43no76zDM05h4qjXDSjdE7o+lKXzj8UA+HbCxXkbzOjdUZXOqHtHDbbi1k0qBsVIo0x9QYyQ
G15bx2NsoyFWddmjQv974a4u9laNznOb0/DmskuHihCKP6ZWfdoQpRggyHQr12WppsEB9I/I0WXm
1wYf4r5N7Xl4uUIi0oPCyc8LsYDGdN7S9ymnz6qJcILklNQxd8VWnzWH6cEp+w4eNTS+3w/Ea1vG
gVeqdN8VjcEzEtMVPJVzuvZvnrMyH3Ogb56qOp1b1Jx4xQY60jdt42zAsmcXGcmSpVYeFTkZPzXb
BvJLoyIszavJ/PBfAR6wR55hVeY8U0WtcfC3jdMKiEhfmKi7ZMZved8UJXQTWWREefPYids336Gl
oe+c9suhS8jpR1EPbE0YfJ3pNxzrx6Vbr5hu2uY2jVrtUWBSGp36ctRzo2TUfW40RIqaGfQAq7h+
FmZMfzZbB6VpIRXoUy8cJtbLOwsH66UozlVdn5UuvJ8aLsOgAs4waVm1IBCtQMx11/JbhoIJh9Od
jzs0+EPFfzV8g0VWffVVc1V+FuI6hk3heLWkrWP3/Y0LtcPkUMIwBQHmaLCvwlVrq0QlooTwv559
HYXBe2tMDpegTFpxg77O7TxxOmf0/Vu1aXjUNwU/HUSmmAuSMca88L1kknnjYnMmIP5myUde+34Y
Yqn0YbuYOZkcGK59tEmuWm3eXGBfRmNJPBpspVSEcFWbvsyMDyIcXMTBoVw6WllhayKtRJrS8qvE
DiSpdfR2Z31E6Ff5DHqsEqfHU7wQn5wIXdzGi2TlSAjJelARss4ZGBnwxjy39y8TxrLqTIS8YUOC
wMzw3pDvtEfsDbJVrKVZbS9Wsi/fkklmU/a60tQp7N6K8dnlJE//ALyQ/SzvcraLUwIWpM1orNOw
jwmcmrhU2ElNhF65ETwDaZA02sFFRYoNHBxKCrhE+riC8Du/wRWbxh/plk13zICFVKpL5DlF7LjQ
gOOP9LPn9x2+bC/c/0hzRva4edXN97scgbbkMdXaq3nwqWypF2/zhbJYV54/Mzkuvw3KLj7GhTn2
zWlcoirj81Ifq60nbyNwh1Ii2uc1C/DXKYqBwJ5zrACwb+zmfJeW3Js6DCarLUJ9fDNslJod4sil
I+VjeSsUn017QrHAMAh31PaeFmKW6mN4sBKg0W51cKwJ9SznyuWULdSj4iunzDCcvC+J2GopeS0T
u5Kce0fuH6scxMuCqmhafE2aLwsAYmTFDZWg4FL10LoDgxeqQTxpLuqC/oMqUHH4FcCgCPhj1rBt
XEZXlcGKLSWVT9AvF9gm2l9ZeAH+I8QEKDWxTalBSgbrKyg8yIGVeOrHADCqdxXrEVvGjjiBlfVZ
SeAZ3jNVRVU31zkfE6uYvGCdV4bK13ap8n/oSdm6QlVEUZegv5zak59rMG91DvU8xozp9EcgUdsb
7RJ4rxPWpnKHZ0tMOwpYKkfsaXjTgjlj6wXVL+N/IUoN0Vlvi95CfWGA/2oADE3gsyWXp7v/x0LY
PAJdtkjtjMlZCBi1Q0b4k1E6wbA1Zts3gHfjALIeAzzs2/91Yy2xK9VDk3peFLaEYDE17oh+SSWM
gHjK3paZs39Sdj2V1UMf7vDS9cvSUkUxjuUyHFThGJqRKMmnGtrnO8Y0vyumYiOOYhWVgbC6IKQV
tODQ3t9zxnkQ46rBj9KvfCkr15H2X8oRrEQx3LSCwxnKF/JR68cmqsdIv8A7tyXBPY7UQhUzY3wK
x0P3U3louReGFnmnkkpq9f8PN+eLFGa+CxDOJXC8yB1sXVqqoBw/ChsDLbRpgv52765rqk88dlqv
C8FMXPG8m6IrulnheuW8dHfgKVCIyTtKTn39bkVzBMUBc4iIhIrthrNDNf7MYa6Vw8MjU47S7SU/
yLh8V0YSskGwzcwW0PrsSlM7u5i9rTH3/D630LfeSYt6EDsmfWMSwqRR532oHQeVxhfoh3oClZ+O
qecouAQXN1bd5YQY1PA8k95tTkCWUyiJMtsUNiCvjV/t/ywmIoAJrF4YyOVuglptDUESJIIxVKtx
sJlnHeI4TGkSVyZnnFxflN8gCNEI8O/EbYNFszNG0VEQkfbmKJ0AMU1BC+WrWKeCNi+bBj8y7lOm
pX1IHLQlEPjbPL7nZdxXMy1JCUAF0q0PxOZtHEU8ftCwc0wCVGEtufIcDd/BTcPuOwZ4gARF/Je3
gVwPnSRe7Vvzk3ocyGSohPSFAJ1hAX7Dj/HmCM+m1ZGLxZ+GrxbJET5IKDIOqELU1yPAAq4CGcpr
bQiUz5FyLhSszVjS8QPRg3pRkBpyEfbl+XANEiYzySGfl9P4LcXgf/XSPDFOFQZSjr2UhoAP5V4l
8EropRrzB5iX0smDKDGoISO5CPqWUMINq5+C5TM3qNS7dpxa1zGnPXvpk9jZgSgudd3FHxbegLq9
acaO6oQSJsLww1FqHaL6dRFDXzfcPZ3lGQXVj6JtkfKj5pvMCwRletPNLP5UQVIF7omXhhE5lcTf
v77rkPS7TEE5IKhpHX+7ho+F8dj1oIenuR+2ISzYRMf7nCn3C73vanLlmeYeu7DcUCyTYA6V+c0n
UhFC2QeyzpbiEzLluQTuxD+5wyQ/eN7JSmvjNLJ8YW5v9YjNFxSQe8qE2bMMrlL1IM/fSe2h2Uni
87mjbVZAkrV4Fcemb7vzfknSTXWX8R3XoiknYwlTG3aShFe+BmFpVTbm+n14eOSTO1UJq5uFQF2D
UKuug1EPogV3FTZjwqn/xbDbno7fj/986QPH8zjrGlzVNN1lns56Hkb7o/svVpEcPUKIJVCZDbbu
JEqtBWrwWdwhScGOEykbdz3uXRvkGj4Suiz1eliWum2YSipW1AuYC/Rz/jZoerS5MDo7oT3TonCp
uOAgUC36cELhy27lAoAskaILQcaG7H/buTUGA5WWsBGThsXwwiM5HUdC5wgMHCH6fOwcnVUZEMIp
smVp7eKdXvn6dVTV96ETbs2rKEztSC6Stm5Pua30y2paKdBZQUzCeVlYbMmKSkH+AeBNWbQ2vT/d
wyHjBG/z1j4VC8hR5IDeRf7ZAFxrRBThqFWcKnnIVLSsen8GbGQ+x1dXwxYFreQQbseqrDWbhYh4
Tx0Q/e/ZeNYTr0gHu9+/ZmGYzQBctKsLyi4fjL1XJ8PHbl0/1fpvVW7AkXqhfSBwjzwrC8voDfZw
qF04e3yF41TsDxf2B9mRzSi9GfLDCH4v51cHrqqNGFtp6Hjh9jn41kJih7f+uSFI+TBkGPxZS8s4
KpAzmgK5Ne1IHDbW+YvnuTjr+AbiNeY4mNiLl+HaIKSaT3eH0iaFc30wbNv03F1hOq5Xbd9veqCQ
RnQ0Zq6/Aa2o50O4xOKPKPSy1MWysYSGGFQOjBciFwJoB1MhI5Si+rdZmtwp3eIyYGAisovQ5jCy
qJpXGCIEv3dnqeMQew+J4iXXYFJVBJaqhFhSmKSsdjivkySuM+1pVcSgtJekpWGbE4R27QfWyiMf
O4Rl7zPDdh3aw/OR1yO7XpEMENJw0NFdsaA0oBO53YomK+H1LREF6iSAMaT3xY5H3Q6Wj7n4FQ/O
1MOACEE+IWM22/d+qf9917LiykaXTEaD1a8GcsbR7AXeFbMHG+aFevRK38vRNkY8tSaXSA16hxpe
N1UOlcqi6SLh5cVoUXVA4DR/qiX3CE0T2UVxi2RKx47L+GkEEiyzMuMwQYclnSt1lkGk/VkY94LM
8C6Z+ERwqyiGb3aU/SUBZfZ/kAdYSBO4XwSqensaOQoZ/jw0MvWcMU5KSgVVTYBTkoC3+JMGCYTG
jGBRNMzRR1V8/XIJWbs2nsyd2A5+dRoN+ZK4ELkXK9btuF3PRacWyKREI+A9N9XeBpaH6e5znPND
VvFjZV0b1lSf1pSimLUc52eW7nRL3hi3dNkzqQC4Q/SooJUn80EqlDQi2YoeS3/0EEOtbJu4DOGP
KEpEztTwSqngGQoYus9BbsSQZMJt8i6iZi2gR5maLS174KXdBWKByfdfCRIiQFPQV3XMWn7PHs7e
3dVgv3VBgE/UCu19+uNUv4/Krrj9VLRHvyD2cQJwHXdkMcX/PAH2x6tI9fvBeWgeFSo2UESxHxvc
VQp21wfnhy79gypcWle4hUvfVXptULj3uyzMstmaAqaTVWRh6avcZWMShuHPnZaO97gBPwNC9ZmE
ZOEGJY5MMTgqAoZBVMaYnq7KK9+fIVzzRq/Ga65/PuP2dGA1qz8YZeI1u15ir+kAQf339PdHOOoL
wiyVfgzM6+pzyk62jQPo+5hEqQjzE2NIUIgiIoQrqX208HoU8CFWBuiOHrebqSICsXeOJmVL0jYm
kjOflVKQwQ190AgXOtDHKoajdDimR3dfhYkDv4E8eHvrSDLl+RKKk9GrW2CfurrXZsX0gIWXNJK5
3CaE930VknySDESqZQzINra7Qe1pv0APMmyEMnBcQpDuuuLRclWHtI2U9A+h0Mx/7fjleO9F/PhG
l5ae7U+taXhrJVGZut9F0dOuCcuDvE+KSU14ffzm41jum1/xR+UpmEe7UTDYwFTYT/uI8WQzqeYi
Dyriq4iLXMT6vFXNMW2K4DQFUsl7Q7byMy7PTn6pt5wn7yUkFYm+7gDepOY4Zks/HOFIqRlUtnP2
8HWCNyzGvh38UF/did+m+a9TyFNMyGxIOaJAMpo0dEe9vvyVSxdyIB/RUFoSRskRPDIHy+dZDetF
xAYZvg9JwYZCLutgfZXFA4Zjov2h3XcUd3/tAhbRhJOmjJdCLC9rVvH8mmNm+bXs5BKN5UTvrv5e
lVk/F8Q4Ec+XRwe8Lo5StJ2yGljTfoXkgSTiiyH4F9XIah8FQdCrd/khMVV+nVQR0Icm6Q5i95PY
E2XplVM4REcqpXcloatAoyeDUTt8sdsaLHDM9GWSbzRjoGJgHCB5Xh+rXdVa4UoiyE0eBlorrirC
A3/oTUnFyWd6TAvBFyWLHrmIThTfN483hGyIDwDO66tR83F9jA+LXxcNzX+Y9f9Sq+Pv2qm/mA4B
YwR8MklBMTEvl3CYLvDqZwIkOtHTg1T6hY2B7uSoSYK0FjWqL2hqR282uNUgCp7sVRHruTK7Z/T+
gRzq5pTpm/Hua5+JqhyWj6zndZnEI+SVGXcFvuuoGr0HjHsKto8YPXtN+EAWHp/cO+EuTadNBeCp
wl/0mcsc+5fMg//ZeVyEKMC3wMQktsc+15arjYHwJGfgLD8AaYvFAh850Tw8p8mvChyZEUgzSIQf
xiKumFw75toHG2C3VktXgc/5Wi5Eux8xFQYJKKyykkcTBJci4E7SQ0NSP2lot2hw2p1LhQUSyLpv
2mAwGoO/bDJDdV038Crp0IpNAQhpTusDS7MjkPeZuocbmBjmGDjoRGevfvgr6pe3QhNkB6hF58a6
mh1eA2SUWvX6C0Fx2GKnENlFpmAuR03isepINGRf9fS8WAwytpzNVl/w2NLFKF6uvVnmWTeocjBl
jhOcMjp+PVq4EA8IE409KweeEBPLrjWVvNrMsg45irNG9Nf7TKTOTYTE99ZYHg+mI+UQHNwpudAv
eJ0XaQNgMf3PbpAm0f6p967bHDxqT9/R4X/itTtc1fn58UToZ6mQIevJQ8rFCjkNARBtzhFcxY6A
qO5PoN5xUZgbnLM+xrikPoVaV8n0IDuDrodhs+WEzbrj2jQ9goW43JL3w+jdCLzHz7HDW5pYUFsO
ZSlCQOueuoSchybwMHLj0/0/cS5BlHGj9mg3+DE5I2aGtO6CwKPDGm26l1SSY9zQFN+udH6aSj+3
83sgGWHR2HjFppHdwSy56ySfj4sPMjfQewHpmW6URAjEdnLPQRs9KdpmOh2Iy1R42F8Nu18NZA8b
krN/U6891J4w4vuafA/IpYje9jgNn5+a+2aCUydnq+F/Zpy197pf8gVti/Dj5Cd+T4IAJjIG9jGp
9sRW+8KT8ivsyriu/TG1KzhnaZOZj7ChO3PqA/gRc8DJreaVW4YDT3OsD7/qkr6H7dVITaACln/0
O73rBuDIRONHT+O5CInX7Vu3tTDKJHJYq2lLILn3t10JLg67shplkSeQa7jGb03Po7Gv6wW9WzFD
ei4tUmZ4DnoimrZ4zeDmm6NXdsE7dr95d6F/8YhU2AeN+Gxb0R/VgYPjFAFxeClH2zSTp8iTB0GY
LB67WR9n+lMbie9C3dGC6eAdYbXhv4OyRnDFok+JsodQJM4D3BFJ0baRkNHnbsJ6l4LB0qlGlMaW
ic9q9Az1v7gXJpDqHZL9TydMmW6mC0j+WBgzlPUc3mXw76SkGzPlHm2NI5K4C3vR8m/OL+oyb96i
+Hh1p8s0lLdalyhHPSJFmCDShUxARsYag4PAf5IeQ5QEi1t5Q72OjXvy3akT5RQnOabofvjY/Frt
gqrfwQhdkM/aTsw1lt/JrZaEhjRNuEJzbhgd5hSXeLKiqtPMphe1vKHlZNW4e0tayJVRobTmQFAv
wZIzU15B57KpZVATZVgL+f8eQM9/shF6ewwa2FIZnAHiHLViB71w5TltLNAsMoJSJepa36oi45FM
LdLTr5KTQ6u5Y0b5su6LwWksMVyelGRmbc9goydqWKovkRi3hiaE35NpRzeEYr9kpleZMGj7J1Iv
B86YRmsHYGArgQIrfkdWsNeyocRH9Dtt4utK63y6zR4n+sXwNVwGBmYKN6M5N81Kh3SgF/+/D486
C6rGX5VhFmFNOvJZj48/Ihrvoo9d+/p5Q6S6HbxUaoZB73b13ZCjPsrWwUaBL35yLKgo1fa+Ygxu
pqKrJju5JR1vxSbVUCTO/S1ls+rF1T/H/x4wZO4kyULBH+L/++QFCz1THoBF+EJeJ0npUzs2wuZu
v5XTVD/8TLQ6rqj+a/4BHTnNpf+YHe+Tq38xFsgwTlXLXP0vrhL+NDKrAfhqTe20ubLvjggjv+G9
EQ+eo3oY/4JYZDCKSAu6xYZ3UEkt1qhEM0D2X99b9XDwXo5GsseuTK+TajV6p5G8iZFU2doOmpl+
JfE+vk2vcAOZ3KcnLu83okhr3Gdf+263ldJx9UzVV9XlLQj0H7qpLzLMkxeJezmtiyHvradZ3qkF
QDH8KNcP3JO5zgzOqbsJDbsh96k25UfMP5TaHdixTA1mIAkFg7v1RJvx7Gx7I3e8ijxJjQeIiIbi
fWGrSktznzKhFTKAmdpfCNWfPgjs8bM/WNpH/iVhS+Xl8eUgdIxvciNsBulbn0TSP0vMr7rRS8eT
D2pq/+DbPr8Map9PWlrltaFVA1vIWB6DT2clAROHX0PPPPTybNQXplpOyKVmVtffnboh5/VLILi7
mdUcgTdp6OPPw9zD82GOKrjS3mAEq4RnTgJdO0m46Ybdgxp6BIlow+ngZZKXBRDvrWZcXQKwFxR5
Km8hlM05lLk+GtfHjOr/xgUzzD9PKxy8RH6DygQZYdsOFncXfDFj6iaugMqcMHmJfXyAuD9DOMG5
OjSVFSFN0+GCW8cfZqPz9pwEiiuhitoFwFZJ/irbkTsg1/AwPn1DU2wAn25Xa8SCvcXueoSt/dsH
QrjWnI4NUn92Pz9iXBl4Zeu18bRETfXazycOZdfwi/KrhdNrqZ20bcuvCINAFxgmSQec1q273AX+
RuvCRHnLf9vTeaGG+Vh2GfhxoT+CHMp/6U5aAPL44WqPa9iMjIlgU6SqThsa3sMk12Say3AeX2TW
7o9SsA4Isq56kQvFP9wPciZxn2wYA0xAZsVgF30pzOeAJdBdBBFt9yZ/5/++ZZGEFcsYuzy7E+Cr
2hhUr/IE3qnZycC7eQ3yOERbEVGD7x1CKAiNzBXSojytv14wI1uPKg8nzlmPNnF3iArqRm4s6NoM
ee3SzZGhWNsZmx46m4jqS4cJFjb13mtHZnmY7rnLrO8m0LzqrvONibUgqkj0pMqBmwafyK+LWpvz
dZEwRRQRbDXPbRIdakLavIM1b7kHlJmVH+/7jEwN6teaBKTgYoE+VX06dCn7Lt1NdkgTXLZDEooj
nOOYllDBx+dfklxbrq/1DLl+XjhhJbOdEdGSlM6t6IO5KDvEEo4CwfUjAS1BAIMjyC+MEA7msb0Z
i10yTIxQgG/cdOW8SthA07cDshdZ7U7km1vihxGlo7mOFIrniOCd2iGOH5Q2zVy+rnQjA16CX5zn
ZqIyocbh7F3H8lBLvsn/6BXLksj4rq8t574Jmtucxmct8pIIvoEnIDnlGVanWLvhUcLCXIVG5g6z
yJOoT5JY5GCQQOBa2CDM0LkUHd+yASNDfLD2C0ZHsH0qjWxl8CZUmpZApra5amCJBGpQhr7da/Yh
oKi/Mbn3P4h+0UO2yldS3zYMGdLDXAsOFhqvNPFWfVqyd5bMmyGsdGUMHT3dtgR7MDiagS0WXxE6
KMgNxTuZ3imF9Uf/IyRyfHGXK445kzYk6FUVpCyHz16nwtnCTzmjQcqbfZeecIIqH+DgPyWvmbV1
b+Y92gArqzTqLHDN3H2j9SbGrSXhMNy52oQrEa+SY2LB7PE7Ax1w2yIT08wY2W6TohLCJV76qymt
AJEdVqstjYUt6WOvbh/3mZkay67IsHAwwVjDsnHyhsJ5GSsFb2hjke3Vv3QKuiFrunDC8KuD7x0W
qQ8nddfF9+TiXFQ0wji0tNWK2tu02/7FywgdLkHQC4AcVrVQINKS2ySv5qSVd7aylWOiU2R0EBFM
gmg+ikT6MgB5CUGR6rcVZch+rq0eA2XCKTiAfVFs7z5btRrtR9QYA0uTRZp5guPBx81JmCqYk8/R
1BRpCMuxyLpLTYJ0IGmyOvPJvFBV6IDLm+uk4JOCNZ4sihrjCSs/vd02gS/ZvsWJrMIj90YT2zC2
AcLSnULO4TQ6NRFpKd/pv3TxDGtnESWU9u9KyETdv1q1oKHLlB/U/Gl/mso+SgafGP9oo82DgD/u
6eTYi/2SiQw3/l+54Fwb9eEYnX8gFVAKmlgprAbjAC3zyQM1IKjQaEtY4eiuc0/3CFaBLCd6D7Nd
xIAd0Rw4YXpfY34IwPvq4oIgBRDl4pLLLTa4rsizQGkdnJjiEzVfuNEzQIX/At9SNuxVcGVDYgRu
bvNUFYGZ+o0rblkVJnCxRYYDTE8oLWuajJ4ylh+kaPkBDXUMPHjjiF+HsHvC6gRwBMKXK8lIJ420
Ymr1khlzw5w4I0cRKDdnOomEt+RBq1WNvDa3tYMEU1OC+74SSgp673pEclWQoeI8gTRGYOj1Rkag
EF+9+mV71dTwWRHYUxM02myRCU71DW2+4+OIyefJ13FajFuxI0c7Xd3Bc7EN2EX+Rwwok7v9fb8F
qhDzUxElNK2ckRsFGvQdEXNM08Rm50wPBAe+7VDqC6VChcxuQJD+lOSpzobzi25eqaYZlYb38XfT
Agxp0/7kgI1CcU8mJrqIZbyvqLmdUUcZPzzrEiWwDgmvunx+xBocDsqVl6+57dLxrrunxy1imeyX
ZFbayUOqoDliovnhQ50iphjVYuJ3VMSKNo/8knO5ZnTHREx3+aIPekCjc8Tn9ZUG/5Q2X/c/Y7/D
R/CW2Q7Yaz0f4mcLgEHW3UUmdHNc5SD47tCHgzcMT2140pqTHeugDV6WZNp8z5Xj8yL+Ecs3ahQp
mABTdaOjPIJ3WvkpQNsCmS1m/uNTM2fJdVZKgphdkPVwU9f8ga9/oDVTCV20veOaQIr9TAWD3PZa
44PUn1i0Zi3z69Sh+kQgXl944d+x1aCeDZXU4l8QvweMk5ttOxhcveLhP8fLZn08zVvYtlXwALxM
39K7BI3fgz0e0piYuWqrEQJa6z0okJ8TLPp56XZ+i9gG+sPZldz+tuq7JzKIzsrVBnA7IhG9vtx7
nsp5JXK8/6q5cFDejN/kxMbwlyzw+XS27QOWEXul/bE+HVCSvSSkIHSzPXJYFCB+HoIDnTWg5qkM
C/YvxsPAUHpPs6nUec/NEO44qqVZBwK8cGUEEHXre1H5/dqq5+OfsulDFazNWJjDrf5/6z1/PTBy
qiQZn2FQ6MH7lAlQVt+2oJIhy+OICCC4mwmMCgnTGFVjdza2uqLo/Fg5qRTDtrl9N9k1j/aagajt
ZfVJWe5wpdyoFPdkOllVMRCgN3PBRi+deOFp861StcKPeoMdekVLbhL6cp/BoqGZCkNnV0vDtf2t
zmRW6PVvFzIfKQFkL4uMbwx5stxaYvkTqtUw4yZpw30JAiQogVLUNY8IATWe1/UA6NubWBFkWweV
a0559d2ShJiXzrCT64ckAbMzl19BntwZsJyGl3wFr6Erxz1kPjgrA79rsZCaUiI9EM1pA7GWkeCO
rwGzHnpuLUZI71yd9OlFhvloOHMQEfzPbXqJECRYguqNSG+I66zVct8HOYntiWj7caycng8GgDN3
9FU0aRBVAIAn2x0lD0z/J95k014G8ZPcBDNvzXubBQcUhrECB45J+/oL0+d+wJYu1MlyYlHdY7/8
VNDQkoX6Os67wqernA4Z6KkIbDh7LREBDGqiGgLtZNlKrw4pNrJ7GBcHY5dwaNud42uipnIITwMi
oqIj5pcFCk+A1j++uJ+HzCUSAdJIsCYQvhFjJR0yJDbpi/1l1ZpGeLFbCg66aCJG+5nHio0Zd75D
Mlj3BITIKRDWE6ZQy1yt53zZUFIBWGMmr1k9P5RXHdEqYiMPchVzcpz7kupBRZrsVcSl0w+fOFub
PRvIksiFimR6/h9h5BYkThl/tP8E1MLlMgNZqR4XnZm+AOPhxJ+f4nYWHF4Utqm4+tsQQ9g37nIZ
QTL6r+yd0nH5UquuxEbo9m1obWWkikPojduLjkwjJ5JoKNSkCKAMSJofEDeGai2zs/13Z+TQZBW/
pj8DEKtLp8Y1b9NroQeH1CIm2TdQ+C4NLPXke6B8SaXFnwl6VK6B7Qm5aBd8rqIaipadAK/HvXhC
4ePON/jeDG+OJ1y7Ir6ikvLc+HdiqfI1pd3wLhDgXjMbgIb+U1c9tHTkfE/jTkkUuHedrr28avk/
n9to/ZLx383RXPkvGJ7A6Z0vDHbSn+PVBeXU0N6576QRkMwuAKqXk1YynuVupTZS96ZMKwuTB9yA
jVaz4VF1bGTvhKsDN0o/qCKfEesnmeGPmEbh89aSkxWjg+VbNk9oLxEK5uKH8hw+oCHfq46MA/J+
3YU16/rUfuMs2VBpOXb3Cp/ijoshoAly47F+ruTgJ8zZBW8mixnPpuEsPEHL/H49u9B1G+g+5ce9
X7p341qZveyk1bR5JREwgkQuLjkt+YS/YZ2PKuXEBxLFEtc1dwz3Oddhu7JpNgeeQx1/nSybOoli
o7dvyaKTBLHYChf9Mf8HpjMEyzyK+vZlJA2fhH4oZy1bvG8nUxK9lVatw4n8XD+tVVkfHNA9IFIy
QY1zck6uYZ+Cff1eeQkLTJl1Pndxl274YQkmvxVdbHXL70WDAT4cXbD7yIUCnmO8We5gak9ohH7p
RHNTB8EmGy7SLoJ8XSZ5Qc54+W/mCxuS6NNjzfNLcTt4TD7Wqf1kTm1YZRIPC8SWbmSutE2/jXHO
UmHMOcWRGdSF4LAlUgWIdQkTI8hS8sL4zbat5ABehptFZ7jcsKeWnIyfXbVUjOxx7dr4slsoh2eH
FUTJ+7jvaSy4cTfWOvnaRuMBD49zeHlrW1Ol99AeG4awFhEdXeBsytjhXSa467ZHEhpCFroCopvm
mtNcJFtaU5ua/ta4hBZml1ncOCTaMbpf9dLPp2qio2Lz4Nnh6upjaVbT01M3CeXTI7/SyqLiVqAT
/MjGVnLFsz9VY+SuVmp/zHWVvpwGu7t70ikiQ1a3uvh97yjJHzRb8If5AC1IqhRWa0cQn4RGskuQ
SXq1Ok13j6icKK2vprDmZsNhlziF5UY+8piXPpOGeM7mroai4hioWnS4ei/r7Q3tHxXYHgr3IFc7
fZt4s1Lfd9r6G55W44z8xTpVtxcmRqMlAkyO6i0g2ue8jHLZ4LkwUki0PLxO5VW0Hf+9wx2O+SIF
rhlGGIA35fLakgGzfC4rGCvUc1kYl310ft2bPdb4DItvjrr27s6pfexzemVlazswKv4xzv9jA+1n
7fMAxvufSmyVAWk9tzPcil2hRpwhdZklxNynPCL9r9wx95a2ifKebdOgW1cexALuJi6upTMQZDvN
qAoBC2Qywzmll1SaC8nDGtqwGgk8UTlddsb5t3oBy1H6Ik+JgyxJZkA8pAGFDeK0+HO/xjqNrdra
xn5/1Y2z41T1wu6LNEsewLCvBLrbsngmG9aFFTh5nAr9fKkmWRpkphj2QxHsmDZ6FsOBvvOQqEmi
h3va98HQ1ysLTM1VD+9eHQXCyU1q6twosUfzqWesjgBHMrPUywe2dWvwITzV2vCy3yxsjI5nOdHz
VHgy4jhy5c836N4l5sufsp1DnJh0sxHCby8wwrW1zDYcgajN6wGPDFNfJceTSYXDFBSjov62AxWv
f+rk8VI7UxOAKnktpLsZKYWZf2QgkPM/IKGOfmaGDKowGXXLl0kZvhEflmtMNm/9mK4wojse7dEv
AqTKFg/2IxqrK8mfJ7cwKoei9byxhykv7pVYdjSNqm3q80eDuFOp2YIpx09qa2TvEPrCzpcOkku8
1xp3iCpBYrU8kSEBVYtLL+dvvwtIFKvPsV3PJj3Io2R1MaEo6XSWqxuxLqSiOhPaL0wTmvFhK1g9
62asc7+s6DR+d9vQLTH0ZMTV7+OmkZdVL1dfzKLD6lKUL19fmGJDPrTbJpzxp5PKO0dyVQ4IiQ/w
4IQtTPIaS8Nnc5Acqx6woYOmCTsPFogJg1gGS4LNWHlfGQkfLABVLcGR2BYHBFgtrtFai91xhpnw
KtBKE8K5Cfjh2Gn8RxWoFsOxnMVzQDju/6b/fk9D4+12Mq2uVUis1Xyu4iSXIouhmOKWBsDqlLdC
G58ygkKxLQu6758sJwnpMwpC94eosn4iuqZrQQz9MrTLOnyqBBZMb47cwtQkqYFu5hTy6iDwPkxo
wXOmkIfuXmZRESvp2TGq8WZnS3mzWaCCwkZxO9rCW1AkfmoQ4GyaWJHTCx/iVdfJy75x6GSjh1uV
Azr+ex37TEquKDLogd0hdJ2G2+KgC7UbCVVtmsxWRzJ86/Gzs621iwAx7oeXqNCTTMyUmde1OSJn
fjYY+q3Di2//OSOwg/aWhT4KceMk1mFe7L5R8ReD/Fs3myQ17n76Z1iAtPfjVGf4YoxWFbOqqQ0P
0ETZC/HHMvCeR7fQRIZY4u+gdaSp3ylHdmYIFq8YJOVBNzudVm4sCjTln1+8PzrirRxJ8v+Imhn8
YUFYPspCV2lTCb7xx0Z0Tz834S82tIuAmWXR9iRqj41fs9Zg/ThvLqiv33hKp6NdN8XtgRBN1LbS
CGVRh3uSK5PJzfX51hHv1snR3GvzeVkkd0To3TSwz5SsmJ/UY4YG9y+O3XHpQYwJCPpTXs3HM7CK
f0gh1RuokfF20cmzZsB3JOiv4rBBY25o7EBCjCJ0kayCunWD6+fk6DfUdl51s5P8mO1hkZVePDNf
DB6UvYUE5WO/8P8YiWKDvdGRtpecpfCSn3Kkkj937wiGspBeKgiJtDV+Yzctb7p6p2iHPx8VUImN
wcSlFeXpCMKFjNGbNkHRJKjKE0hz48yVr6rV91SImjr1JyVG9UViFeRLvzjRlPYFm0JP5Z9639S2
RDnN8YJwGG4zSAryoujzclV++NeCwCEWya7QFuw2cQN3oYU6HeNq9KoEL5wbS60GcnE9r41aODOg
K1ZVqleFGGl5mORMtzR1PAxt5iWZfT3qitaHKEme//BcnvwP7NG9dkkguC7v3JA4fz7TAHaqQWSG
JlC06SrL0BT3OYH3hnMxAp90AC0FnvKQErR/T7QmBS1/4GeXBsyN11oGjWwZ8HhpiC8Crtp0Pt4h
5w4ESXljljk5IYDISDA0mU/JDLuwwqAEC92wMvZAhasqCYiPkHxqLyB50FBS2MUID2WfEBiqBWLQ
Hu8G4hMhpT6rIcZcKQ1jKKsKIzQqeynPB0eBq4dIm9dIBuxXLUCN6tEFymTLMzGKEnNZmZXoMFzV
OwE1WsvZ3yPc88Cmz40HYHwsmheU5oS6Yq8dp1Qw+P0+GIe1AuG/f3gXXWAAf2qZFbHybJQTy8j5
XvpS9TNdWq17nG0N1UQcx9QyzIKXbhbj/bVuWr/KAUrUzrA0kTRDcuc0eaFq2PcNYmNOQFyzQfMv
6jnqKQWeBKDrY6sRpfsqusI4/p8dd5O7OHoO7mIyG/TfgH1XNt/+L1O/JkeMACdAOAKL/S2/RL3h
Z5cujKk2Dt3/wj3/JtZCfLZFIC7kRjigBhq+xa9QneyoCqB0wtzampiiT5EASrFEElcaAsbpscsz
OWmlOaE1B4Dtgl/y/X7eIOLXbyGeM/SppVZHqwLs0J18GreWJWn7Lteb4FOrtdfJOpN1q//AGiSw
mtJMgTIasK7ke+LsuDmR60/oce+MQjPh+Vd14g9WEYKrzTNjbzbh6XHhJDhHYy0cqlcgnds9MBLH
X/c6guiI/UgfdkBhNY3gdATkJ0Bmk3wcr5slH1ByKUpmgrv/YFYGAWS+qNWi+B/psdjnLbAgqOJe
2/oX5wYAY38sgHIg36u9ta2iQnFP468nGYj8XgCSmSrEkX8/IDXmIBN7f3aX5GsYsExSqSlnkTqz
f3JKSoKfJC/cSDrqK7A6vjJi5uhbsmTwhE2gHTwXdMk6LTb3fNNW1XgeStvkoGWecKVFymDZE7QG
Rp4ajfQWamL/R1HJzR0ifeXToLB5zhCzEBM92QDFPM1jicWOUZgx/7shM0XwHDptc6BMf33FI+nU
HntbPL+GElizmw2if0glKn24Tyo6/ucslhKs3dxI3+ik2/J/kOPy9Sh2Y7BnWLfgyLZWbUldlbSW
bNjASN6YFZ+X9ip8XqEjKr5NUnMdMCLMfs4bbVQgOUpXCbvFhdvkZfO6iAyUgYm1xDs2LSocoZto
lp8f1iGrzSvumHCjEq+7T+dU2Ef8IUVNvDnHvunbAFV5Mhv32IhD/Gosy8Hy4k7w56DP2FUu19qH
rtT0ORIYXk9oZRRpVBihm7vcx0mEPSWceFLeEl6zOYNa4WIXRC1dwdL1P+YEmIp/IVzxwCh3XsJm
tXkFqOzmAPk7S46JinkfEO26R62+AbouLZ4TbNkxcbCKQRaQ+mTWzlxsAJUlBGpOlNdpZkpBPIaa
vxKwG13DfZjYSRQDIkolEtOZjuj2oLTBG1Kkm42h6bE+ZoU/KyDuOcnpY6naJa3ITEFyeGm7HYAJ
IwVkAeu8+wrICmbEpH+HRNhoeenKCkf541zSnXNe4YY57Sgrjz33shKGbSfevJXuMJT4zTEQ1O93
agZub5tI3gKwUPsRcPnzWbPN/eOyPUCU35/H5+HMFGF8UJZK16YcIHLAzez3KxolfMg7R93YRFRf
V5YuXZbYIe8RJMLDdzRGLFNJnAy3IXmj3nrkr0Vk6SqD+XcXt0D1N5DFTs7jn13+34Tp1oQSiiQM
0drAAQ0AbcPaJpKumxynPsVT8O6KGWTMvjtjuPiOoBTZX7UoeEiliwaE0X3RUvEAfBuBBMAQmd9L
I+d2zvbtrK+k8ev71BoLbjCOu6drBF3KwE7LAoL5ljZQw6Oh+d+ZigEgQQvZT4xf8x5ioIpbFueW
tqPKxtIccsQirLmX1utHdsHOFgv1yCJHZjZChTrpIFqJF08FmU+o3o7cVKs2TOixE7BmH0GkOv0L
L9GQNFw9Xa+zml+Mw00yltVo0T3SRaMJtO5hONCAPSFS6q1cUcEoCASl5vO+0kN22ukRNXXnSdrL
8EeheTTPNc3bX+ATaz++E84UMC1NHSWEDLPl8xiEMiCmSDvd5v8cuZNi0hFv4+KA0oIh5/cbHwzo
Od2KziAdtyYjePrnWbPPKyofbT3RQFxbpnEKd7/niUpvhEK9HefJ116X5CXoB+ADxhKuichW60hU
j01XFp8zK786KKah+U3zOzGtcSSAP2NVz/lT9/ET+/fvs/zE92+z/Z888ZbURTZkzltWTLQcDeVp
i5QmR9JXH17pXd78Niy55iDJDiqs0HIbQUM8wmXFAox6sQxXOih1SlPUz5pzpBXpezVDi0tu+cyV
gX6DnUzvprtvCmTLQEGflXziYU5RHH5ozW/p/pBfB6K4IKxIn0f6qKAbh1Yv3vNNlinkGxuIMJ6j
ASEf0LaJA5OBXevKG4x6m7mP6KDSbbZ8irClQ9JkAVU3p+7gVFRnEnTyR2DbcBUq/xMoO8B9eNYs
qkU0ht6QdGLCiqQvFAm1AlQG8NrPipwDH6bGnZChJWZ6coVFIAV1S/wuSxZfIgBMoKApelYJdAly
ZRKywkBv1E2AtQXo3gLatfUbjXmaR7m0xP4ZPMPK06pkg5Mqcyz+n2d6wGHIR4S7ETdk2ZRFNuTQ
yYEx64JhHbxIhfXwhoy25es/LSbXXXOEBD89t2VdjIGnGeqAJZksZz+0YFDOowFQ+wjPaDzf9Kio
/nieMP90RvM9SIxTl1451EjqxCDLTK2YtnPXXMyfUUOGM2JFoiyrjYSv7jURHHs8Ws3bMPyN8VMt
htpOVI+NfH+r1xEaca9BXoPFD8kFddXo77+F/S/T4z7wd2LiiZO4cj/9TLPsx3cBOH7XxqmpKXp4
ZlMKA1QLFXw+L9EmBDSUurI04zT9JyUyye7sSfASnU1pNiJuxkbZOUSDFzwcvvepAkwqYoAyZE59
gZV/pccfC6a48HYhpzgGVR+AAkwS9iDvmobRfETXQaNdXTlfFwU3gTbm4BmNfky8JorE3bogEDob
k3xUSXMHcHJs8DdMi1wRp1BkkfoGUa+EskNBPkxLHvF/2qoUhIxA9Siw8vgSpS+qvloQLP5m37Z7
0tYfEFYPH6jnfy/cyHTF9OnlFfEaNFChkBihWV5k2h005spvKKwwk6UIt2NjmqxQrZ7EhTkqnngq
JuxKYyyjSCRqB0ojLeu4u6Td1ScoxpUou8HX8c7TLcQFvR333qbK1ZntlDWQbd6jxRLAre2StEfp
PnHt+L7xMz/fy2l01H0hWedC/rkfPpyoTZtsfSEbMSFbCP6/NLHU2xjPRYuf9YB8MNKfENp4j8Wj
oxRbW2rEcJkuSqjsOg95B8d8iPspydV1F1mywtRZpLDDOdeYuRMz1ckGhQw0GNAmh48mokzmRsad
p7ajtRQP9IrGUFy9FkwGy4PmALGXoRDuFVtrY3TPBk6plZIYBF8Ob9UbcQEO02aF/69OX2Pe/5vh
Fl3xgDj2KyRKu+sZ5w1QbDeQ8yCEB7LpcvWrqninx6Se4uKsv6iwm+qIDgBLFVMJLLWC+i0b+gKj
aOBDgx/ejG3t/SOzO9BqioyXEaAqGzrDa0e6U/dXDVRi6/GaqSjA+FR0tIVyUQCpyAuYn1NuUkQa
j+izxZZFkYsVM9Pe58Hbe/5IeaYjXU/nyJkRF+iGFQnrilZJmim7qfvrdtMKSvWzFc0iMPreA4jH
M/yiJkGP+2Zc9iwAeDz6tEz52C43fD3gYheWDdBkaP/RBBtI/0OtPnxmyDkQRdd4f60xkUA8IFZJ
zQ/qOoaYhidg46Q7zb4gAwgTiM0EjkJVIUL2qxyjF9MPU3c2RIi2GkzprEjIv8KMx5jm7BiqWx3s
xU8haCZDpx1a0KABaip5SL+Zfa5cTKXUFHNhMBmwNOMNsPwVYz+6XCOGrbn5vZmmSudYBrV42SWj
chZmuxV49Y/HbdmHKTGxVRii90kIS8RiGXzC5foWKlyexJ3Xhd8gyhWgBhmINQMKiL6n0yua4Mr+
I5kmXyE+6cnBq8L0zGXZg0eLpoFf8OYBYOQkGHMxIVPzMyXZ8+uihm2r+PGiQ9F1fPfV6LUMB9bT
mFuv+RmPQ+d1UjqNbq0sdi0MOnULo35G58ExHCSLONdEDCdVHndp2Pjceh+1JLoPu49vM4PM0AFm
10/fuG+P6VKnXkv2ayqDx730bprAVA3PkzI0rNUejPSA7izBpI3cBWrzOHugcpbTZsR7GEBmQ+zg
m+GorKUv8r2oa9j7ya4zavryIb+FIVjsSTC0e2BzIatDTUtpIw82JM7Be/+nkZQOMzIdPuykCKHF
qhZCKuzjv1ejXCHQz16RwsR8iOLYT/tHN/B5V+wc03/xMggVLKjCLCbXI47C6i3REp57OdNC6C89
tLvvOS8SIjo72uE/+jIFQAzHrXCea+lf6UrrPTysL/iieS3nirL/eULIAeFzw78PN5J37AkYpRGF
jxRj4YEufK0BLsDBbnxoFDWUzX4waeNx/1yuhcKrEq/0BHAWcKO8u8Tvu4ofypzgEQ8UlXT7nr2E
m6GhiOPtHo/CW+zE6A76X5KKlinytBMWxxI+otK1tzUS1i5qkuDN1jpLZ0k3F/gZkgwtV6E1ViJ6
vyH7p9wbS9/mglPXZFRmcJDMieU4IJfVxJEeUujJn74Op796DPqsYQmz8W71RsQWiinmcObtgKH1
lb0nTd77qmwLzt5w7qm4vrycuhRKWbe9RRNDWooUmMecqj+kgdMfktPlCn0YZv5OJZbD+G+oogjF
DYkeyPsy6T4eTwEa6DqX2marcV24AJ4XF3qVnGzJPEderMgKL64cD89wmvck5Tb6U9U8eQTqBiOm
T+gc4zF6uzr0RGCKkN/nV/MkdJuk+6KitJmKEl8IEmNXQpQZ9YKXjs9WIXQE4Wg3fU1k9sB+Xh9r
UNPDpnddUljA84eqDLDbd6Hu+5W6uN1saPBG3yTlXvVBT9VafuSVpu37ms8I+O2sjPJHFYe4CZna
EK3A3q9XiL0Z0r8VoqIBbzA+lagxAi0XytmkNEzVJMy9yXzpv4JcGmthLIks3iYmjzGVnef5sxXp
1mcG+KcR4LAa1J52ktP+BOzXNdmiz+r6r4ZG3Pv1K5S2aU7alREjvxIXtalC1AixX3pH+x8xTJpm
/qR7o5/0CJo7ZJDJguLjqzPTQA+0Hvkm76s3bgQVK/wWKn5MOaKlDjomWDQsWaXRhOUun1S7z1/C
5JQncgTXnj3iLGRCfwjqg4cKEpCvovl4bpk42l1112mOc4eHiPKMxGKILbBZs0iy4LKl8DtsVnGz
DzO87Xedd4vRU3V81BCLhGX85/bcxGVX7+iQJpLe9JshjxOXP74torkeQ+tNhSv4+EdCrJEXj2FT
MpoRPcLsx2cgK9fsiDOVwaRgJkN9JXseCGiLcT72jTPewlNdmC2BLiJj4iEeeUaAI+3TwpWuYYWn
XdNeSu8Kc0DiIC5OcTxgwq2fkeqzjqJFjPgVZXntAFbYOZg0AI5d8lHdnvGqxiNr7E4p0RjC+5Yp
OQ2OgUumO1G0sAHwu7DmRdFDImIqQ7zGwGqAgoZXWHXFxKGaI3LoVk+XIst8lkhm7KqurZh0lxPt
vOEF/AoCbfxRp7aRg2f75/010EqW5O6mmxcNEw4XQCiOCvPOEtmAgDrAKBdA2q0CO+TJt0KMvW2b
4IyPmtF2uska4AUZ6RCcPe4qJXve3bJu9Bwgpn4BgGtzOv/1vWjoIrvOefcPAeFPpg5nfCF+pk7G
RJoGzXCJNZZ026EeW8bA+dVXfe9sW6njDmPFZbZnuVO451QhJeTleBOwTFOsyWLsyPBnUWvi9YSY
fR/rRCM59dX0JK13/dCDBhue7dit41zPLD9DT5XyyvIUt9weZQwwhWy9U+qWVmtwzRouP7XwRf1i
bBCnrzF6kp5aQe6UCgjqRmqN853pfirmg5E+UvnQGc4NwcaVP09kWKsIQ4Y/FqwCriXN7qNQua+0
b1T7f6jCkT2NZYZw0GKg7OWn4KelLUkP1Sr/mk+LVlGGNEJQaaw+TLjdSBiI5OqILgI11Gt/cXD2
MEAs0l6WDElSMx1ZUcmU8hO/cU36GBDYgJMVV8jbWlwdHSvnOV5ZtJrPYkucKixE5N37unIuz7Tj
j1kaQefGCWX3fWdVtN6SHPt8ZRJHe8sFDu9xiycDC5FEg+UAicwhLjUvTZTPHgCgi//P6YyRb/yB
suTG792pKQZoIgayi8fuxkcsp2g0ykoAMOu3LUxTS4GoJ4S5bbtHmmHcz3nuEYoGOiYUwV6SxXfC
be+xKR5Evs7Ps9B+PHKmkrBV3Nkfb2UwnpSGU6jaZHjvA3MZfvqJFmAVA7EOf+8rK6UfpOAQIRAF
JpPPDxXyUmGp/IVjWlmHzpQoOcRxP9YkECXDMtmVH8Yw20DXusurs66YR8TBqjGQ6Cku3mJ5k2Mu
FiOdtDuFjks1/zXIaYHwf19q2a1bFNPbBLxKZveLSMGDDdD782jTuVWa0rPHARaK/VW8Smy4FWwx
FDjhGhG9+2V4q62L6rtOgoiktLTHrsdrSXI9jyNAN/n8Wy+6a0jHsAtXxe9VH/ZDd3ZbS74onaha
5QfQIyyzO3y96MamDE8xjL6eLFbU0vkef1c4ojnq8/9CshN5ApMJ0xnBJ+T/6sdIc81HM+OI1rgz
l+kibXvX5gjOinJ8+49eQEk3hClvQKXwDsjaBfhjlfTFtr9iEFDGYOSCg9eexPB6wExX4wqWnD5c
UjURwbwnWS/yfnr5LKoaF6JiNV3aRtyF+AVjlZPLexUtWXNWQJKtJ7O3c34xysLcN06flJD1LIX8
Yf5ggHsUWgMYuHTMtbj275fhdGVeFSBrA86n6sN9dSdCEK8UCshQ9iu4j6V9X5juzvKjTFLOYYdS
rlJU2Z9YubTXyDbco97ub3E7w4KFfaf4JqmrGJjX/+f3F/RdB2iXfBg1fOy7sqc5tvB2sY1lv4qE
UirJdiUwENNsDuQoO6YVWxMESuYVrHtK7kWglK49kpJt0ArxL3lHXUyD4Qig2WE1+Yilm6AUXtAT
PA2nfnPP8SlPEjKdNr6sLaxKZX+jacpgP5EGB8rnI5rqdaToV6jgkG2a6pJxcMZVSMAWYOIcBErW
2KVqoft0Wj1k+0b9uXTzpIoxhFLGSM/IEBtgXAIKkMbNqiWW2fOpYqSjrxCiEKDmnMIom7ovU1NO
9hZOHWqks5RQfykFzpjTxtM8xEq1hAj/qbQUxyS1W53+/iM9CtUyslRmK99RgDdS7VBqBGoaek7W
vq892IMW2dmNIOt+ymXLYHUQz1A1jJZmzwUNRRXktL84wLu2sadPX3MKstaygYuXS1XoOyguh9bi
P4dVro0sdDFlR3FGM0eLJlDEQMWXniNNq7X0DHBSmZlryBacJH0Ig+7t2YdUSb8bhA6x1vtXggEB
jZdbg8ljNSAx1RKAfiz7bLaSJ5mwuReaj5toUH1oFXwbiShxueWR6MbMZP7dQAMIWWm6R0avDtc5
L8nPYvYfC4wPjaDibXK+W9vcr8+zZZpq+RNJGb2GjZi3LHE9PzzoAlQXPVGxb2/8KLJ0QsuGjzSd
jFCosPRgE5ATm6IBGvSH0mJkeUUbONhy5rAZ8NWjKFak3hrb8LmP8SjDskaJhil343wgicxPJgEh
gzwSV+eYoCgXIis/bx7t25xhefa6ZJGsCQ4mN7fdEiYWyX6MkXEFXGszA4Brbrt4NyfjW8m/pKfl
g4YU06iIdFiI0YwrPOpFbjJbZuQw5a9dabQX4Wo4WU12NJ4ZHpdetcHH5K4w4dXNdnO+7PD7HsdC
6hVa5BCMLZ/6Z1MTfwwi0rC2GzNOeqyOttzekKYrtsaz9l1ajfbNkZEHmsfpW8vkvlLNJdniKQKe
f5RxCZeAjzbAAfQwvGYxgZYiFKa08zU85D58U1UhAFS3U4KkYnnlTReFOkAdA+8QnmwlS+7btXkI
LBfqar0hdmjIzVcYFvO9Ft0De4Y072B8jqod+st27i00Jbot/QX7QTwiTAYGbUtSjTfZY9S86Xy8
hwehzD8KZC0NwZwoLRqYuFJL+G4hVKHhx4aDjkzQBfE9gzGJJiPeNwEBlnGoKwZgotJ4LxXXjVll
nkJWU+Qxg1KwvXHdpKQ/W1wEb4ofOlxw3ZZjyqo1AD6KXhYQ6p2F3COqH2yD15NHfiLSil4w7KUB
VZppipJTRTKS+D3zY5NW89Sa0nLL6gvOeo+EveBOMgR3B5H20Dy0gDHI0UcuFB5kOIhM5fWZ7TZS
HDovk1VmOZ+2+WCpOCU4KJbp0wfJT4nw1/EprJyeeVzmVVkJQ2giZ4ehCi688LOsW7NC66RQYzAo
1RwOEQwK/B4PBRF0ISQ7Xys6tLNWdoJWzmqakdeGnmiGKveJrgsbDrvrRC762j8uqGOktn2RKMiy
m5FQyQPnvb3hm5Z3IMEmB4b+7VjyuueMZwkE1kdZE05cuTixEmh1GUBlA2RBHgKlHPawZFH8HuXd
VHGz3IjozBG16S40hKT8t+8/tfOucPdGmBRvlXD1YM0IUW9el1nQK+w6mNlSBTWVTOzZEkbecKP5
am7pLkl9CI/F0UlMrJTBgMkOyHk+iMgCHYGLlNg8V4W8WN+sQcFcxGkikq+H75WqFtgwemBpO0bF
7b+BIs5JK4DcGGXdRyHCna4fTL7f1oZNLGpXgPQNjvJGiulJ4eGlfx05J1R5+Mt3xDl/q9ngJVmc
QCCOL7aKwsobdvTUDiw8Dpu1W6cFrIyOP1W3ce0VBuEe68ScoFlenpX04FXrJRxxwSmRZqaGbuLN
FCW/Np+4B61WDboqqvR15933zDKC2wIPwlalAFXLWxrPK0wZt8pU+pgr6JudvINQfgz5jCc4bMO0
Mr6wh2bkWy0fMF1p8Bn7I4F+fJTaX+M4N/8Wk1IT62r8cR1E3/yGuNi3VCK+MuBs92RIiB63I1Q0
8s4GEA3T4SJ1EUuWGEoHTlvxmKscdxO0jy9+gIGjNyQ9XQx6/FfIAriZ1tC3mUcGbOiNpUWlIjOd
6eL15nVQksP6dJNItvD1QFjNQ7QNlRPKk5M7pzfKO3V8dyQRkMQU/sBIMqIFgfHdEGYxFXy2uV5x
mr2rBqaNwRQdahxRsTcxGPvrLvca3QOo4pWPrN0JQN6GAWu5amKgukUBnATuoiSdkDy6HBpDrkdn
N2pif1wQ79PYZpi3/IHZcHudrR7hg0rLssS9GQCLQWMThzswE+h+FcBWKt7CZXImZqAlDmEHtwOT
i5+rVc+GE9FH+D5hJlrJ7b8rTaCWjAjiCgjN0OzjPzUKSovd9vJ933fDCAWYQ9oYEAVCqV08m71R
nLqMeQsCLaKqHO9Aq+a6XTLeIQcAmc+dO1TJyr+On64nknbVBg5ybCfiP2sziclFoE/Q2pgg/BOT
7yUEE2+MA8XT6A3lDbgVRWIInUDr5Pl0ILEuq1U7bkEl2JNied66I13mJ3vGJS/PgO6W1hqFeASJ
jJ3+S3N+FVZcV7QFVbtv3yUOM/StwHdV2LYjbyIfJuo5j4ZloDZtXZx6ttSVPn8PjEGjgUpk80/I
UjOFVcmCKxQgHPlJLfB+D58t8uNV+3hdgJDDIHCuZNEE+GippbxNMYHpSdlu/fX/FW1d3AGze2p4
keFwS67jqL2xvXKG6O/uk/FsZ2mglRYNB9Dpk9/W6LoJWVE0ymBRbq8gLBnPKwtavcgGtknvhQCM
4pf4D5J+VKMeobYentxXkfu5+olak0dY00ZENZKCiVhYvf+Gy6+L7IN1W5c+gzz4M+8cDo0qauac
daYdna0+graK+VgzPrWVzj/UDpLKxme5k1/8MKpfKuBMIuI7lfWZnlOYV5MamMXlU5Jantr4ZKpM
X4WdJU4eIrIqXHXCCfaLcYBb/Jhvbsnw3fYtz1TBng4tnPxVn27lLmHabVt+430D4QZULUWGhlOa
KGc7h/rvMutSUgf+oFQbuBCeADyi+utwoP8r6e/JeCxRvYOjjI6HoMJKHzAtv0SaJI7fr3zhfqqX
/OBF2+BSu62+sH6ya30aGvch4ZrfW8MMXU1/y62nHejJkQF1WwupPMTVkOGz6aacTfMq50e5UUwR
NxxKvUa/bSCWF+dvHeNPlSm517jqsd/cR6ldC5xFHKHoLOp+DfbQVACoYtsKvnO00VRBVXgdvf0E
591dV6GT/nU5/euHjttC/PKB7KcEs+y9/qptLlZ809t0JyHScT6UBQ3KlpxHr60mU6KRZKPlAehg
CrFT2gY+DBo/5kK+Zpn6Vt6cwuG5MyFyKXihqBLo6pIZQCjvv32hKSQHvlfiQyg+N9ZrtOw+IfYi
1oZ5apfcL1SSOJCuKe4WwFh0vuhNRMuEwR8P2LT1FIg8pBkziKoFYimKIcjHDhIdVr/YogBg4r+C
xpWRfH9kjtRkHJz5pvM6oA9HzCV/7KVMRATHy/zQict3YOAzQXS/+mu8E5f0W9ETN4TkzlE7ytIh
Ey72UqRJdYaTUN04TtZHGGNpmAEdbRXsYvEFQyUDaWOoQsyHcs/GJ5TsKTbTX5ln0gRtDfI9aOhg
LZjC2xbLc2IGSSwwdkWTmLmawzlTwRD1NB+KSr2Dkm7B+B6kYwfk5T7pPjp+oWld/npGeXm5sJDw
oI/nBYzBY3NuQFrl6Z/9Pt8b3UiZs6vZ0FRYTMAv3L2b/ZMVggBOe5lTuBml+1sZFoY7aDYpndva
DGEhu7HL2Za6fWsmh4/qqi3AXjSbc7QsB7RkvS0tCa1XKukpJyXQ0yaU5wqPJ3aUd85T9bEG0331
XwHgkQvV/ieEF6/Vl0rU3LyPydQllj8uNg7a5TxD7SFzN8ZL5NR3PS2jRrnAzTl3KdU4tV4Fz5MU
UW/Rsh0sDdImDNBmNRkWIB8cIJoVcFP0bZNJrVnryDIVtEMlYNvmHXnSNIZAwlWzL+T6GZQUzH8L
zujM4wTeM64oPYMSksySQogt7TxcxHHRtncnpMWfBK59Y/Kz1IFS8JdXlcLUvEFKs1dKqUsnL+66
DiIQcRgFGZ2YvW4bMpEHW24tbguxYWf3Mb9hHDxmhFHKu0sT313mTCMTUS4+h/I5oWyMwu2LXbPn
dCvBv3D/9xhsfoyb7kY2k2GrA5zmEgsCUEiIbHkS8jsUm1wcSjqwt1MZgwwELachW+YqsO/V1tUl
j22QRIkMQiJkl07HM9y+JBCy6VzrcygfMyEPDPEEpwUSM8rCIF+c7/OOMZgOiZ2XP5b1uCur3zcG
F0EdL5q9nFKxA1ZdD3zUJSoJFLSOK4r9iNwO96qc5mEzfG/UJwCX5mtwhr2V/r6onmDdPttsXSeu
UVlJ/dQ9Bt1BUUwFud8gudfBIscrSZSDx8FjGx/K74yahcFlcrsrvzaqDM021dQ2304Qx/CRUwPe
QImAsdc52kLcylx2pOlYeHDPbWhFY4rCaymsJFW6G60YMGjp/iRNTf0QLcd92bGZdUgIBium8jsf
DA58FW3TeKmpMDseH6/6YucPvlI6FfA/6zZaThSs/YfAQW96keeNy/wxhkr8he5+nMOYA97oYeq9
x58DJdOEeREuGf5wpBvmLnEV3mG34EZpfgsAYAhstriU/HAQ3bS/mBK7NIbYrjmoQJ/iffB48Dzg
qpKPswFxCgu7ALSq4QKK5M2MLOt0KzqsV/XZDeJiSGckD8qH0TJH4d6/+1wQiKZFQAc7uujJAJoX
9oEJ6pO08ERyOXUMdm1pz2eo3hZAL8gkqEe4kAWx07x5A3TdnUGkdlLW3JYMAtn2pKASTwEfwflt
+2mUN4dVOPJ3ucPAAzs35HlkZ8kWcKeZhDnUNcIXjcACyXtxbE3TbUT/jAndnV9W/SH6O5HvU+0V
wzZcmyDgwkibJAxWWImoIzrgo/jS+1iyENlFE9Y+ZOMSZXNWusAOGpWCNsTl7bEQlbAFkoH/Pu3R
34lmcqvZZnKRBf8tkNsnpCFRunikwT/c/x11g+oC83xAzs7vYxs7od7qBaivMxui65j5oe7H+8aJ
+EbzW2c/GYz3nzAXsrX6o17JRg/sJpi0Vac8faQ4jxLNLmllUBjdpPSwEUMzYuwYQuH1jw2LJaJ9
hvD9JwDBJ0N9tFYs3l1BYnwVVRTNfm0JjG/d8TSvm31FxrswPytjFPbfVwlcAiBzCBIsT6A11kPA
rJcpUlz6oXFTC+0d3gARzFRef17WQKGd+HfNNR4WJ6gzaW0GdLEZotXOjr/BpuGrVEZWDiX3ROA7
LQuAmUHVmIwHd3Pze5cg2i5inn5/6mij0Lv5J0zbuu1F2YtdAFKZQsK8/o+Re8h7ovUkiFVm6x+o
V3Baui/qHkuYsujYWCmA9K1CoBVJJgVtfmW9g4nLOF8nFqsMC6yT0P8+Qlmpr+5RwSZhCvsiuT+V
JVC+P0ibAf2H9Y2+ALotiIAI5nnxQVhIx9CoJ85ITiO+QRH7l5DO+3AecbemhN7Sue785/De4KpZ
GwQ88kDfc9Y3GMAnCdnoNiOUsXiMoHyFUeosx1wBCTmMzidMX0mf1TAoCHAMvGZ5NYaPhpPldEeC
fIQQ+YUI9tUivCUvlPEP0QMBTBgH5621UDsaytU25vrQqD9UlD8Ch4FcbTDBK0Rxx5TcXTDYw0ia
nkh9l1ThZ1NcqcPKaptrXQ2w89u9gD1WgpO4ZZEZmVUfWuO0hGn7l5x4fowe3mvgoF7T5pPMT4FA
YgGB8a2Aa/EKmJRQVPHTkrpeQ7H0lxf4Tvr5VN5N63ZvNoiUVobDlHnLdGtnitbkxp6a0HrolFhU
Jlq87IiEz9lflmIZbhlK/X+SEXxeOQJzq9e5QacC9VWXn/K2atuFBmkVF9DsEja4/9yzMpPY6G3T
SVya8Q5IBAaT+/7pyrcVacmXIoDBDP3jEx+eEVgIkPkkq0yJiymlvIMoaBDbmjtkMCo0L8Kc6+YK
XUjNFrLo8S8lhdIovhHrQ0mgiin61Qz11K+Brl31UHxwh+J8ylBNMxNxTV2KNhk2/cu2mhNU9JYT
JaXX8j+KxcsAzY1QZzeFZ1vYKr/NHcjGncs4JWXSiulnWU3UESmzMGzEpaqB0lc52z3+uwshO9wu
ZOoDl0P/lwu2FY0GJh1Xi5T7zUao4OEMRGEeadtR0VisF6gGhspLFc1+rhVlKJM+fzpqvDpiY4F+
uGhZP7uzl5cv0ZWvd2XNINU9M2ZHtGkwrE0v7ZJZwS44loyS356HRyxH8GuBbHupRH1crvnq+ytR
1R/iHFQYBPH5IUSME6eoARtYv8QyGzSXAk+zPG0u0dnn06kR9oeGLIRAE2fbof4rexCaPvHRWNMS
isJL+NBe7wiNu49Q0bbn5Y9gIkaVSvAzRChPQL3xPkc84Us70/bncusVjsQfInFiraN1vAvHe+m7
T7Kr7i65TL5I+IqXD4FMOuZ6PqfLkFFgC5j94e4Ov/8fMsySwdScOmsQxbJJ9SxcFRd/fw07trOl
DWAUP8LRi8m711roiMP9bbVzt6r0yc66FWe3+cKpglNtsOPR56jnsHNrOTG1rVohUoNdz/12OhZx
1mXipReIir6SyI91hX9nvSXqZbWl4HoP+W1tDmCo7GF/HIRy+4mCEVyDaws/rWnHQpCWX3stMlwq
xlda8rw2CCSquRcfHhqlZo3B8hQKORk/ci/qevsidbGLFFAq1cTT/xQdFnMcvc7kpqzIQRi4XdIT
7B65I7l0wHVsDdXYX2DKwTSFZ7qNzNOUIg5jI/UMGWHK74RcbSjQz4mQDEpj2YIUKTCgiPB5kePF
RLz7QbkONDR+LnA7+0EdhwcOZSCL/UZ4JCpFwW3nfoROL5IzqxCzAmSHprNt9vhYMds5W8LOiUik
81seNYCPNmq6xyySQ+Ta/ZDj27H1t3p/fGlxECkz5Qh0QkDOdTwLOKHACeQQJEpw1ywAPoiZqJ3V
7TO3mYEgjxiwwhAK8wEa2EO61d3QrxyN1a2wKmSN9sNyFH4Y8DZKv9q/bpDoh69c6oXbOi/dDFOU
AcZSL+o6G+rqyRGsF0LRkFP70GEzcNeEIXOYJuz0I2MJYLPvnrajPEMz86e73Y3lYaTntPlyIwWi
alGk05FXS78PiErmDxmKdGxQ8EhxbUu358HpMOjAqGHJuf0Q3LaYB0u5w3HCYeK1EyAUEV1uWcGw
Cv265Xag19EgdXTSZ1KhxcLJaWqAU4PDPxRQGRrKcsh3OfezHpKS+ZaeweREab7iqQxG19yqVuAh
/C9EvwFnLvQk6oe1HjhCkYCUFZvXgmCjHGjHEwq/eNb+hh3LkYIobHHrRI3Cv2sjXifEj5O0jk8z
AJl78YYX1y0DCFIWkdSlWd/XnkvBJtHtC7oHbYNWZ+2NBfgFIMok5G8dbsJztKy5D39MqTFyloqI
c0dKe8RTTjEu1ZI21wWuI0Dnw9iBQuv7nlLUqzKfgPoqOJJc4ogSQJWh48yImITcJO/V0BlJLIMR
RLrbkLyx+Ir5pwkLnKrP6py2fJbzY9sFmYXs8yWfQ9kcR2sBXNAb+N1gszyO3YJlrukoMIjv+xS6
FpDmMja4Z20wWw4qIqFHLLgCUWiobNLhakZlQ90FeNPvErKet9HCsb/Y7HkieNY2B3ddAAy6AQfG
vYgK3rJFoQybHa4Ad745ZJ/mCPeyFfktlkG0Kt0OrwdJ1Fqg4b3UQTgqbrvSsSssT7oxM8pVHTOL
0jEAspAQhoyLFzC3P+t3SLnvjfcoEgZo1+kfBXyK78e0yAJzRctVmaUZfaKqW/tgvjq/TG0rEHJe
0iDlKzkXDZonE0QxXvYGzMc8a1L2/L4EHCiHsmVObaoWD4Ghxm70Ig+AZBZWe4IZdOMKmyaZFREG
+/mCwlsw93SIqdhrsBjMSs/YtGkhCXc6stVorWbavZxq2V0xrT6a7nfjZy9UMWTembXzKnTkhKBj
Nknbg435tPbATxohV6nLq3u7IJ1xTKxa1fCDTcZY7FVCjcdY7E8B1UJV0X59DHDmy90vfdSNf/3t
+Jj2AuYrFNFWBQ210wGjKbXHxbngoI/YHG7rCnUBDOkyg5+SeEVoG/Nr9hlg4VOxCdDZoGmZefDK
pSSlqG/tcXzERZhB5cqdZpI3CZREFKEoOZZez0cyDbj9/x0Hm8kLqsJQrIgLnvPHRjirqHQ3F54+
gDakeQj9ho3b/oIQK2lcwPTHqZI5ANvStg9gU53McPl581LUEySH1lbZaYPdYyvjmHSj4iSLynsN
U6Rk4EQ4PRNo9dHNSxD8VBVN7btaPGVNRTQUBiG22BJ7QS6R5K60WgkVR7zNJ1A2l2J8WVeZt/8K
6SrYA01GGdS8maD1FZbdj5OjozeUaZLcm1LaK8lVlyT/Y6cFJc8BngrxuBZ4CZNp+e53zCWfmVcx
Dz/Rp1GmEZHT3of10tKxRB8qmOKekrrChIqka6FQky6okeZtann917gAc6HR7O4naJF0NP4kxEVH
1+5gKXR5ANzPnzFT2kOUXmlA9JjAXOKNH2kq4jpfiV4yEHlBni1gY1rjSHqLCiVE5gcBgV9EAt0N
banp5lbjYg71t30SvHc6FdH2wmgcHZwNS4bIHOQZx9e9Dj6juCTqbT1hagZPwitLEw7JuCD5CdQY
SfI+0oNmySpPmLYvKnwoNPyiCgXFi02m2ECJeXJzjc/aZ80xeYeTF2KfXXh4ElbZAZDMpJqEUvXP
5cPs45zi753C5gLOEFviRN/h3mKp2bcu4voxaSiFBj3kOlOldD/iY9OaDZ5DTvxA7ns/1j52qUho
P60GWcQgaxc8IA/QPuLF0F0g7mAy8nG94vTcT3qL/0+lf6zbm+roHas26JI4HqbAeKHP4Xzp7kPU
WTiaM2mYtR+cjCM/rMIrdOHhuQskZgIHQE/4qrNTsiVhS4C6LlfPy6/wI8R69pHOOWmFoloD8a3e
wfqnwOMMOvTzsIu2FuB2mopXr17dO6ABRBTf2zRTP8Vh69cMc/DSp3mBThyVke+zTWYpyCTzuXnA
ENpywynEPQRB9MCY1+8nUir5OvowPyCJDZ8WD/lAteANaBrsdU8U+J7AYOAv5PRDWUjBmF6zlaQZ
GW4l6YJP5dOTlhk1tmBuDZA8eFb42sFIEObZoOexo0UARk68Yxm1yPOqJc6gXOQAJobDklzAXQIr
+2PiOiODB9Qa14YMLtKZx2c9818oodzd9FJsosBfCs6BPk33TkaOz/0RT+qHuIzKw3nkg++zjRgD
Tbz17FjY430kz3HzFOfVrkcUDezpDCe3cr38NWk46caBEonhCpZ+aaoiBc+OkHuAY9BZuh5kD4sk
eZBXHUkSa5l6THhsHXk7l9OXXzmPJ3BgZJ0QNDGKuQ7xwsdO6TOB+MNt/5awKLEQp6sXXF5BqTtG
QmrdV30mwLdwX0M+QlSTI7Ta9MTRvLC+LS8/GqTw8SdKJj1/0DW/qIxfdVqav/G2qV07s9aZEJWG
CEnXckNURonONWAOjr+cawjdLhTzeWdB5Mj639l4N1qudebapxuCT4hW/YVPyUiLp/H+5OT6jFNv
Z/zClmKOA5hzwfVY9QB29Vtpng0gQBk+vEgteP8ZgdqmJGuKE0741E4gypx0INN+26UbgNd/QIR7
SG2zSYh/3UdorKeQf1btjh04j78QEJMVzkmRFsIwL3Bc+Eb79etuLsoFQJTsBCL+dcnmHrY/hGfI
qT5wR3BLEHXlOGaCsioboplIMWDy+ivoq4AWaj1DeDR8s/Lnt396SGzMJpPGpyfU24+4Mev6obuH
Y1iyYtpAbp7XAi0+9063ajaB3paKW+exEVAl6s+/H7JNTLUIZ+mwl5evUW5EG+p4XcVEP5w77S+l
sGInKxtJdiwd/p+BGJXRHJ4wCw/i9SDBQweowAawBwyRpbiqNitdbwMtqaTUumccrZ7hv90lVkjI
EJ6AAD+sumUY9D3mUtNRqb4SkzzgpyQPY9DSRzfTDwOFT9c5HxaX498HllPYjwJQUuPpgkcSNS0r
36p4sbeaq27QMCSFQXgWukVUTO7ut7vHo1HkBdPGTFB6Zl3unh7Lq0foDvQCYUlam6QiuHsdBvJi
VNDEPKOBBCjKHZqW2fzeEyhbYE2fJza4g0jCUoY55nZY1G/4bmhc3H9x2zgPOSvCQ2FCwiw4rPYY
JsJYZRfgiEun5se0TjmqJYFoLhktGcy6cOcd0Vt7VqkMEQBEiLK1GpuqtF0dBxdP9P/msGLJqOjM
qFxHvkU/XO+dtmBmPXQk/DLBBs2LP8crs3oClKW6/Vu02VzXeW0RZADej1zD7TaKAd1yxyL/kmxU
5tRqeA/XwPP86eGDIw4ZaKdrIy00gUe2L2I2l+pS+mABcshNJF5zfgGElMuo8ot61Sktvi7EItk+
V9moSs4O7uIYyyc9OUOjMdqpMBxWqnvG5KdOmmKJrCmHYwE5GQ+KKp/YhuduMVL9cGyNTXDEdKcA
gA5Pgo/ENS/DTccIuIPsehmUrBcwlIOWAGB0sUEFZty/MttczU8dgu6sEOBuUxFcqWDj6JSs1hpv
NTUNTPR97q4OoYrMzvcTyxCh3qZwmitravmnpM3ZCedGQ9MHWZ/tuTorCHMWixUGegIjIRc6xkc3
wNrXi8TgKSodybdOJzZ7x36cg/MdUcqb/i8v0pbox+q4cmINLN9OSdQ7YWvcBBvdxO7G1hUqUdHO
HAdQZxNIzXQZzRiBsZwnG76zqbca/QP7Rv87yBzxM7J1KUY4bbIOBB4k/c/oXdSxYJdRYA17us4w
3O8TqkF887vYt7HH4R5id6DZjTxJBx/qMo8+VGHwCnTwAyDwOhZhJnWgUFkS67pZBH5A4aY20VS6
6+xRDGpzFPBeuVOwF7wrq6EWbdYrjl9MSmqSBH0GrurYB0hmJL/64iDCKf6qmpJ0GKsn/aQPbdcc
DRA33jdUi1ypPBoxWCNQOpEAFqNeGnaCZjo8Q2O4AB1S5qUW24iZhRG3nrTnYQCCjQH9PIgDvCSN
7IzN3JyHVSdecOtN/ibLxTOys/ROVBuJiaOd+ZpSDcWdnm+xBCSERFb/zAWN7aZl1N8040+3A0u7
HjIVfIjVlXZ4Uu7Ca0dRg7s9v6bWlAK8qIboylohn1Q8bb+muwvyKSFMFH/LzAgTkTNKUHuESou2
xEWe/jG4uxNJusU2j/6vm/d0Kyc4K7fQp91JcWDSxs0Qdc5qL+hppTIyxZ/ZDM75gKUrDrfebOUU
aaS9TWOUavyU1rjBCtxh8HNNVWleGDmJLtrkjoo3espuWowI+gUNpfxjg+zAYVwXeYtrSQpo7whK
YVwGZBjJucB92aGGW0jzTcVGP1etFkrc4q924hMwkQHXcybTNUDJAHuKQVXgBr9bo2xaE/DEG7kw
5S2Sx9Bb9HFDZgZfCE7EWq6TbE48J0Y4w8cL5w5jRAanD/S8bsADFQsLQxYeI5gWRWScsIyiRXo1
cu1ZkIuzt4k0Z3GI/mxJVnnqyJdT+3nUL4VCOnPDYWkWsneLsT3WBfra1Tbr1BL7ZveklpDKg1Am
c38lKtY1pjVNLyS3Jw1mq/LWKM8EGfguKPpc1x8e2PpOLpi5w68x9jnY0GEuEt8doreO8IARtOsB
A3Oe+r18dzmiY1KY3cju1EyptG6OlaID8kcpPeUKjU1eRIc73vk64Yn6IgapaNSgrqW4GELmyR3C
FlY2wGjI9iqme5aBX0Y5BTU+s9G6TMLRt3vsVXuVLq1ehd20GFloc2RqakABvJ3n2eKuIqokr/8Z
ZhTKDW3cCIuuix+gkR3xfLurf5HqVggZ3GIG9cE/1utmISE5eobmoLnha0DY/Dimr+CbpQvq+Brb
h2aIv7tN1ISAgqZipobR0mIdn1C0uz46HusOh6HgjPnyiGLraUBgydrQvllzscQUkC/avh0YI5j8
2/YnVv7JnbDSKJcBFhQjSaruPDFqiWabnq2G/jN3ALJBxWvg5idF65AVPu1dOixAwliICrIMi4Lg
Gw81GUyTjVyv6tc3OVB5QBG2lmvV5vmPmQVlq2fs+YvK6pHuv/5ng+PSykdKevE3MsyW5e0DjjkN
6iCLKuAVlgLngUb4BBGlqmQBexaBCEHaDfAGKRi+lClltzUzZzL46kZZzEQlCkaWOoQNAY8eiktp
3qT/PK24Nh0oez7tAHRvVAbhFaQ46v6hONvRcL1JBR5kaYVTWDQol85CepXt5LVipVlBK9ftwhG3
aoWg6jBFaJWhAt75fP4PX4GMTtFLNLwiuyhkP+wEGcxKHp7g9FWqABCm/ZHzV59BJCPAaRPtPFFK
NO98U4PZEM+BZsoZug07/WzlFIEJVMMH3oHyDJQNnkb9SJLwcLvFhpl8L7A3jweB8Kz3+p5wuxVQ
WdzPN49HXyMT5xdPqMHG+ODgUcEQ4z5fvuo/pQOk0xrNh2Ztuu/W2BKjeMDYgn4PSvTb69uu6Z4v
AiEZhTwr/RkSlKPtX51Ulw9JuqWsIsgkw2ZcqlStEHuSo7E9LagRH9aamRxnTWMhVBEVdWqPTMyE
gs5GgOvGKVfS0Dp1BY0q6E3d/Od8GK32yWQAESMUUrzt47vOLQailBRGCdz7B22AzcYowIUOMyAU
YA4/nmQByDy856RlgBqJakUzvtVUlx8oxb8OUX9QaaP0w00VLHzCl2WzS1mjap75fV/ghltAMe5W
mja9ZleFYvpYW7luOAdftcoOxYxYCZdU6NF/eYBKYmM2ZsWNPb5SHcb1cCTbZ7LtSqpiMN+3Rlys
ji4umogbnKP8GNu5rS8sc4ZoCg2N2kKk4vg9Q0scMut4KXWHYNaWEU3jCUZ0rAT3xj2DuqN0jnhg
4449HP63TgIBMrt7hU83LS3BSJkIDKl5FXEs3UlNK2bGeL1tDFyFNpSlQCcQHuU5zQM1qvDM7Rj+
66ClX8syHXeM1T4IUNevaJNzFY8A4UOf0xKaqwOtjezBYzR5dHuVipCbhAyValDBaAf1n6sFpyxR
eNmnPvKLcUYsSO2a3tc9mRG2U6sme6FykGzp2N0LVrk2+/WPvE4KC5bQYN1DepXzYmTppERHlbIV
bswyP1neJxFq4164YVWssCd/HWjI4M+GUmxMGLktwmo3hL1TkU0JMQYO5oVCmcFv6oALXKQcQvTO
jnp4ZSc8jNaa643DWG4qb5t9f9PvT6I68N0zb8cV4h9PFekezzI/eCPhDyRjAmtqWFbEN3X9pnAl
z0ojD/9MZXhq7tEStOse/SJstFU8UBTyZfZV3qlezzf1R9WsdJntDRwl4DGJwrTh6NvqOKiFpYsm
NGBIgXBk5fI7SKM06+YEA1rDc49IWmOvqur4veVUHE1AcmB1rSYhDuv6pMpTKPThTEt4xHZCqh5v
CARwbElLvlcCMZw0sCYzmPpmxajEcln+ZyJ/7i9jTT64M8jcFX3+l6qnyycGyVfBxBYin5JktAzY
aEl8lQPpYeHrWbpiwIJT4vVU3n5MDWqvMO5dbyfqaKCGeIrjWUdq9C2BVpEZfBC1mH9EylvBl5cr
a8sxjMNgnUcP0EtPam8fIxRd8rVTclLRrSr+CQtOsnmjRAQtewtQ9bqHV731apWvOg/+yJlQO2zn
FPiUmNmqvIBg3mJrJXXD7xpdQB91q9U8oKqYAUIsiQhfEYeMxWuFR3PlJ7IE9hrkru05JBWGv90x
z7j08ihhpbbsdfol28JAvLVpRumhPo3Zs2gmBjT8ARBiU/nQzhrFxBzcJr0WcyvjsV8iM3Bsjk03
Y6wtd8MeZuHn0veKV7UaPFb5tD3fA8rZk8dI1hRHO6+uSz8VZjAsqjnltbFm6JFA5ntu3GyZjKAC
ydDWh6pAjsP+yfS1LBhZZ73fqDwou7L5zql3d2CKD+STY5s56gxm1TTAnWxQsfJrXTepMZ84iscr
4WzNocPdQKt4szx2lYDgR0JHpElUDGLO7kFY97GkQyrYu+M8qFZDIKeRkmdvdyjGLut6ShluSfBH
565FMCp/1/dJff4oz5ob5VTH6SkBcsz9nD3AQNz+4RslYltM0Jd72cXUM0aDBk/ebkLhInnKWHqJ
EfH0zuku0K+wER2JIbt04DTbKOy4lwrQfV7tv7vwaVYOdGjyPO6CLd9MMlw08CQy5dd7OBIJWDNm
CzN02G0NgRrlyduu7+uWVlflN8o4kBpaRV+w7xvwP0dSYHerXnDAIs7hCsvE0FAmdoT6kjs8B84/
SwHh779kMfLPIRdGSOWuGT+heWm/PuFujBdx954e1VadwoyqB5tghbDm3Ra6MqWsJPfmUexHqTgh
ySPYT8mM3BPHKzP+OEyHiwNetgnmgwJtnBa25KdNs2WAiLJmtR7dlh4+WA/idiCZtC1zonQ7subA
eQBY1/XUTcQ2RPcgN8gAhFjHvmnji/gc+wjfIoh+5zGN2R+CyVjF+58vE+UqpdL5/TDXbsGKNkD3
scM3RbeEqOjA28UHsvOeMqVvSbinaSuz6Uh8Wt8h4bg0ZbgeptUXr4epzviw9C8Az8spS6c2MCdU
3cHiA7hIFi6S3UdNxkKYTO353IX7tyAVlMmFibPPit2nrC5W51MLc64KQCuqpib9aJyko5OWIz5G
ZCbJVSj44T/E56n/o1T3q2K75nNp4R9OlrH0OWkrBojqf073zvJaXxcYKZdNWXAmm2CSoyWjzIGn
xhwGm/uDLnPKw9GrzWV1PbP0x6NK/ypEUNv2SfYc6hxT4S0W+qOudIU7m1nr4mfHYQ/5QY3gub1z
Vem/cIUs8KeA1MUseD0sgJqJz04E4koXm7mr2RUIPN+G19PvykJUKKCbHMbcsUCIyCyTC4+bnpYF
c6gTLKP7+s6PNdKo4KJzposGSE43k01h0YinrU1oswA7rg3dvvGwDQkjhK3WLldTNjQPE+PmcJ9b
huf1wUyibQ2a54oOzrK0ooEpOkvXUE+/G9wrxZ0KFasRvKzGk6Joc9v4V2M6EhFwaeioSZHXGa2Y
B0yta5dRHMrcl3RkgAk1aMMhFHulKEpuYyoGmfWtXwbgitNAKmM1P52KlxoWTFcxmBZLSLsTY0G5
Z7+YsXWYY+XhYCm8hiF4W56HO6aGV9CchS/KjFCPbgHWAs73QvbWoH3U13yZwbKv9sU/J4f76A5s
MgxqcUHuxH809Cuyl2Kk6W1IBSWQjvzw6/enMbUQ5sq1P6hG8HlY9ykbG7ieNdnd86vOQH7homG0
O8tM96Fx3uraulvN6zjOFhboOL3QVIEXCXLVuNXfl1RcnQqCtdUkmTJ5myUapJHQ34selITyeOeV
VwkchjWz2y6zew2nOzaQ9r7sx8ChK3sBgUgbgsZuvlKz0G6kVXiXeECrybm+jw/7RDCi0t/A7HG7
BybD7wOlRvT7V0HiwTsrEn1684Jxe6hgqQjgnpDdXl8Y1Dp9U8oCDTyjOqMOmcRttuuxxrIrrPHO
YPm7DlnTIM9ajHt5N0wAmZOIGT41iHReHMjw9f3bt+WwL349WRjILp9HnEnidlALG1ojJUGnins2
IXOLe50UqZkxrYqWaRbzrAc7Rgkh/G+oai64iAZ9HsnaiGvoom2kviMGroVTuIPaxnbUX/I7jjyW
IWjZoNQAOTvsvnrJdxFR7Ej46AIWubwJ1DQlyXDAARZzWMsttbpjFhC1BDVdJAv8LD+1Lxdd+jGL
312tY5HsymfNZHHnIaGuScj4pArtM2o8QFYRpl6tOLBCEDGf7Byptz65hjzalicFOWmoygfqo6N1
W+ktuf9XNVJsV1xv14o+HoGsZ4llHB0UPU0hHvjXGw6W4w1zzVqSknL8/wd+1zMlWMhVvHe1WnBg
jTePhFa3nlTjpZlB6hk9pnL7S4veotkjZFAA+PllhAPBQf0jLnlrcJbiKeBWrhDUK4wQjdRJAAfZ
7SOOgWngXfZ8AFuZffpvfR1r/Umwj4whosCP6O5ffQgiV3/w1NoMrVZnbDjtxr8TT1Kl3vkQ0TKl
dtWppTdYh0A652oPyK6OOXgU4P+0wC4cDrspaN2MCPX4zLsB0e0WeBeE+08llkcwC9yw+nxMsW6k
zXFOo/0ISo2tKZc7bRkJTnBOGCg2r2OImQ17ozSCWZ8Ej/TbxBvcql8pH4uyNBAtIadLvdkl3aoA
dQoujuUw+R4DpFbbB7hnOSGyIPRsgufn9ZxiLeTal6dYh6vV3aLs82R7uNSn6Tox46fBLus+65f9
2sFGky0OPWOEySp1FoBEyAGImyeG3KpGA41NslXwJg21bObgBUUwdv5uNhCpjthoVhroOREsnwMZ
htqqWl4f8qRSMP1+EPppKGaJsUqN6Wr6OXDBmtRVPJzeRRbm1tamEkttHWXhHyqRAUkpnFdyH24g
NNmgbhRl/H9M3x9DmZL0vGdcA29uThfNj5i+2SHA1AAutZt0E7VrzBSKOq2qH0BkZ7Hul7K/pUzz
+kaBVXDqbEZxBBP8Wj2UTCbrwRYVjH4GY9wqZORE0gNDuBNWTkYDjC9QR5oMfLnCVctEgR51k8dw
1p5mKdM6xG4OZFNbBfK6rTaGOYO9SEi2j867e8I+da2vEngF6bU0TJIz9ElrQraSNE7tRnj1ljrh
MOwt4koH4VKzmrdpAxjTQyNFzz5DdnPhqte4qEgfa3OtcUkNWKWUHcTPhklmAw8Dx0j1wNOCFuHr
2Qc46svHZmuXq5sVdDmPmgaeThMOWIn5MraHjT1BD/X6jX21lrVzG8QnXeVvd3Uj60xTwKoGtOzb
ZlyVcY/4iZcpQA+3O0QkbOKvZPwKWxEYQyso6bkaIQCpHxPT0qiRLwEhHL1L8ll9GjH4xhPtVvez
OuHLzP5UgpiKfQ7dofwP951v3enPqQn2gtqH/xWP4+4H/eOcXR88DLpugI/PUUIGlTV6EbirA/ma
tPeDYUr2yG6fhzexusVtG6bxaIcmmuQ2Ztb41jxxsy5/hYKrwMWtgWV8sRJi8Nx4JBM4A8p0Ajzc
m1+8yohMUgjxnP2aQ9m9ldQop9Xb6RGMxmirz1B2nPTzSgTqOmtRL0g3TkFGEEVDVmnUvFf2HgGH
S4RTVnxPQEAVw5MdQYkVmcqqpGXwY5bRm+WhWAUZktB0AEWq6c2mk7KcC/ou3sY+SRzE6eSoH+Nw
MDIVUP8w21unTSMqLK0LDwJzg9DGpSHQr15zAYef2AdTFetZG9G7B2DiBUdyvs8fR9cOfhIx7O7C
QBVN+gB+wHuV2e4n0lDro3tMFo+O71XPSsq5EmfncVnjjetOG1ehnop3E8t+40A8S7KwP+MTEh2R
NOMpl6LqsYiSdoPqdcyXTHb+kZbekqc2JbC44K+soUUvqpS+Qx7A9A09o22WmKcnmc9jgHLZMjxZ
zKbOGaDGNXsrAk8SKlye50Yr5/JoB2t52K8DHHDq3LpaXt7f/RZG6UwZRXX476iTWi6iQf6E76U6
rAsE6maHCQw0aiOJ9dEuXfd9HbzuerIZ3p+RhM9zNjBZO5pNMe+txyQ1a5zYT017PDWobCkbMjCG
qB2v5tNx+F0JGYjqzrVJpTnCi0y6lagoBj7WoBefDJdg5kBaZcJDH0abUe5heEtbMBQrqlyuLTTd
tikFhf2H6yue0N9zfxA6W9Q0/R+SYECTygt8A2SD9XgAcfNJNL2dnY+UgVdSvwk/1Jh1Fx2veCyj
1IEmbABTJ4tfU9JP9wjN3ZpkvaI0ivUz2pPmulMxZ639S3nFYRNeO7FrWagQ3SvTWHi0XJKl15vB
kZLTeDmucDTlYdaEFd11PkaHxrEKH+dJNLH7vKqVAoGYzaXklsZDuKMbfXgWb4/IJ5FVDc6AFc+1
SU++BvldvvIvNU18r+poX6QBCRUgtoNTNUIo6+ndO11zkPTuuWsmCj8LjqDLzXtomI0gUBvVxMIe
SmACY55U0laW7pATkODHMQqELhQ4ZiaYbpax1Q+tHZ83B2lSFUtFRxqTp9Wz6urXGIRTydaRooWR
iCG63LSlvrI80gkwrzrbTXzU7UcPhZiFH3wbVPNTJGbSRm2ccqdH7bmyCPsz3Fn+po+z/xVwswy9
s2za4P+RoZOKD7xlFN4DwwkGlgEq2QxAxHPPGP7zgygPh1SqCbbVJ7PKrHTal6H0dGA8sYqmjtQI
mX0F2L7s2yrVViFdjG6mpZF23IbU999ZZvIuPMhOiY4+7KxrcjC26f/eire/8o6GUFfALy1rnG2f
0izenMsedQ3gD0bkjlW5sw/Juua3de5ON7drPtXqBVcg1ZJSZybXZa3jsZGes6/vFGge8KBCUPEO
WVJ5D6w5YRjjRyQ33CBYIq329l4HRcM2UdcZoaEQ0M908FD6DvWUHYSFGPFczpceI3zb9M7SpjHG
qSii6EQ/SHyjUzaqpzJqJMsyeAMBG35eB+8wFEu+tY02FWY8Ay/wDO6TQSns/lIbS97WMFMCPh77
IRHpHlnlr620VOd2XnsYxAIFtzHPNxt6eptjP4UIFMSxmBWgDvdsSoZfe7g2P1UjK1ghv9z8pgl1
5CqMkDaCD+XgU5AXosbBN+iOpLnxIJlmGM970XoV3UZ0BcDGiveZ7d9GtrD6unD5VCx7OjmSyLaT
fFNRCdZSf6e1Aqr2ofcdR43J1sKz1C3GHviYgOVpXnB1QK2386VPfFlemsLwz3yhAClHydqqPSuc
kV2l8BRzt92rJLZMsa36C8QsoCZdJd5NqkuK39HYF7U4+KGvk6wPEbWhZorye57GPsbzSWw6D8EB
PbNurENWlp2/a9RSIhvnMmk1W9kEgiGWXscwjBCPCzwggveoWmJlsVduzgB/b5V4MgSMI/kG4s9G
N3NtzXWteMBWFAFE+bB3nciq190kcZoNUsqDsbTYRRqy5yWOlAdwklJcQIEOzUiBVq5QMfak7Yzl
PCG3LzVxEw7NOTLWIsV66Dy4kGCVKug5uY+zH4ytbBHQbXx6q2SBih9jFbNtqx8bGEp/MRUthi9r
JXIvVpMrjCZuSAl61xkPWpGlEX+/bJDX+seFm/evzazkJqOo20jFlr/Hia9HqNif5BxSLTotufNb
6nIyCAsXA9e2RhZiUq/nJk+oMhEHF6uC55jjA5H65QA6lTq9xjyL060ZVmlG9mhbf1imSrBd53Yn
GvSgyvtVupSxYSYu4otnbY2N3KTZC4jSMmZIOB9c1Q0kUrxDJw8Xq4JYYFZWrvq4KVtaUYtzzFLs
WgWeu73l9S5zAudV2pa56A71+cl2BysTzicpYUwVC6ovrG9wn9CVFDezPKGIB3gaXloERO3pZ42A
LN9oEpv0ADQW1J9dOjzIVq4wxCHrA04xlkwS6r+IfA9yQF1qHxONO25JU3+hvzNxO/FXgbD48gUf
ox1r2MWXvIKx2LR1ABlf9ahL5EKkeZsU/w//LZCHi1+zAB120ERfe1gTM9NCwBH4BRXaH5BWjF1N
O5M6D/Glw7U/zOYZq0kZiyoL6lMrWQphR9fStJSHE/pT8GdDcCodun1s7f210CF+ir31bMvYuLA5
kKRDAuGf1aZkQ+X/2Z9JGeVxdz8/pYtzasa/cgVhlWryO/9D6WAMieISR8U1n7K3Ude2NwX2fZue
MnXhqdxcakxiKUQE7lHjeExdN7UXSFakSOBNkTKdDj+ot6lp7BNcpdgKM1K0FHpoInxOAe/Y7xDt
baGI2DFZ+sBvoBwp1sVzA4n8Maq/rq6BO6+hJoOCO1nTfUJlkif1GNQyISAsBfdYKhbdK8+zCRjk
De/syvP+q435izo2aZ48RuaV7uuOGZS+Q05+gQbB+Ad57WuJj7QGw/sk2whmvEhNbMDyuMpqWHVK
yfyGogd0PMlmto0DN/683l0lmJc08eHJkC0Ud2YRrzD6wkCs9iXkHuGAu/2OlklrBJLTPCTGdwcR
pABLBHLWV9TcsckxhiAJCSqGHy4/GEt6tqPnNu4LXHQIWuWbHbTlpMjcMoSORW0qoyTUS4wQePNV
zdGfemm9JxnTocfAeuHeack5VSn/E6/fPpeWq7UMmUeR5qo789DmrM/5/pwz/ZCiZOIqyXUX75Bc
ctuuHdQvGxrgHUrVd7h+6tBt6xgOVyiGMO+k+gpdxnDvOZjyTAbjRnsP9N62CD9h+Udj4G4Xc9yp
MxEWsYeBkGsdnPps//6ak2n7jPZVXwmCQM1OooM7LI+kaRAm+ggHiQUJuwjRRiO8lKco8IZGRq0Z
udlNgFBNCedbJhabkVyTft93qdIG+AMh/AIIXLCVjKIgb07haamRj+uShZhpDupDcfo23a/NUXfX
bGa7WwBVtS+smEclR9duSlOrAbIMU2B1+tA605hSeCmxU2UaZ6iTf46w1vEQZ28/yuUxuOEWTMKL
l3XdIahhBMuCAwz42ffiXE8XX+SYanOPwq1JnYeAjZOhEeQMCoHklrDiSKMqCwfbCrp8gCdHmLtA
XtjwgTuzZu2JxTm8m7rz8ilVzQU15HEIAWYruKrqS8oFsCBR1VIGmZsAExKTn7EtGoCy/7Xk/WGu
UDa1lj35eG9LsQANEWfC60QRPXe57PFG8Birdhgb7TiiTi7s/6Hx0LLcOEAzHHOMrZyizsjlcBJv
lvizzO/tyMEUfmmyy5KsReeXJT6hKvIfETNX5qS/wPIWzFRJtIkhOjujr8jJjGAeHjJ9EPXieLv0
h6U0Auc4jJabOKR/8nFCXYkP4WiGcrypeOHtq873P71BC4/c9g6ePu42IFTqLczjLx3TA0gD7JOi
fEL90Osnk0ngnY3KoYWgmIMSRzMGNiJ5Z3ROFUr0agr8yxkIPRIT66YwEIMYPVQrfKWgubFkAnmh
W/YBCbU+D8A+Q1KRGJL08RLG0wEv0whi2GGfUxQW77fx2pRDJAqIfKZrl6A9eFpK1nAcx8tDUq/5
cDME9mWfvjbTiq//ZDUM2DaNFBs/nresL3+syGAWYBg1b049YsZnsR+Usts3R5k1drW4UVoWGT06
3wag8VXO8syxQpW7z2S9RP0ls8e4YyNyJa3r9713Bt0sg/3GiFUdiRgNADS+G+X5W6F23fvsCpgP
93jKzNfIa3ACqjPv072dGfttaK5xEENY20kKE1MY3Yd3tyf0Q5aeCT5YXHsF4xrMew0toAtN0Xel
SWcq49nI7E/OO/iEgb1Q81prdKg4jrsvZ6rf6BTCy/LiCsvFaJkfuD0gXn5eoKvkb9AtiuhDC7Ug
ln/glKmSDtncG3aRiPYBpN5ByJEczy1wJ6FyVOXXadCEDLVXLLv7Ba7Gy7Omy+7sndruwLFrZXh5
3E07eTIHexTMssVfzhiIkFjrhjatjoRJflMBmihq9f1Ll/Iojd38IfqSF5zRXWwJqBnCD8hWfQLV
d4pTVV57P2zPB9OVTPUu+bKdACfVWtqErCZ9qZZgNpUjEnkpgJAnRzZiZM0lJNtciCt/P5SuO4KV
m3SFYWkMl4F2N16ZTcaGS7gpSHPA1JxktLseems0b/ooTQBw7BckCrvrl7mnBTnErbIUQyupN7KI
5vcWjhtQ6qax16V46Ayu74mjOlf3rsqv7AT4JxrcXE8pf/7z12UxWwsb7wnkN+Z9H6kaucR4UgmU
BOomgF7LQ6JADDm33knKfwFxU0fzzIFJ3AlHDsWwn3hoAOAmygSyywv18VkMbMw7TzkNQ4IHdNWR
/D8mpWqba5WBFhfDRDi0MC0YsdBdIcsCKEa9bjbV1jLsYhsU/WaruOUQkxfrmLZLBanC5QFgpD5B
96ufJ9R2dd5YLxmaPCReyjiWjU7zolo8IoaTLnIXCDHAnikHHMyvP/3QGLo3H1Aohz9/Zk3xaPGp
Qg9zGp+QpX7ytWUZAEdJTF8v9htMeINnfKivMQa/LpzYyGH3Wty4a0azVpPu8UyGcr2b4AN/wFIS
cfpKjDiA0EOstkvM8Q/lPJXMq5ReKNXjlNs6eJ3V0rpXrLxp31Fe3Fx0aCvFwEJj1PPF7VcfeHyL
E1NIRln94nN+gYSj1XwdbWNf0NNL8DscWOcGHyOXOMF4F7sFIv0bSSt19w1U0UqJsgg6hy8bBHFm
4QElyNUYGnFDQE8BcxsYI0VZD/UWOru4ebehxPr3icUoNGIQ3prN2w6QDuae8c71BzfhzZew9Az/
2Jaq0JtRCjL+LbuwLAS+gdECkq9TjAl/v51wzZJKUEOlt4f+MlD2/ydg2e9LN51TwC3zljDzn41/
DBOrQthC8MmN/DCn11E3q3dGG42yvf1cRqDK9gD/ebZoujAxZ72WqnS0BP7blvYMgs1rl3+BRASg
dolxXr1usVsNZs/LyUPswp0adrmEUFLaJu9mcQVTGU1nrV3O+ZFb+12yL6+Zlll/ldPg8SaAPPIB
8HuSv6cWz6Wj3RDXSaVm9S82OpoUNkoCy2Fufzct84ZlswVbLzJEGuvLyKYjEr/2gROuxZ/G3Thi
VXTTsecQblED4bUf2yabb59r8EsTcjhNWTR5YR1BEwDuq2eHv1uUTSnZV6D1G63mvXrLQayBoXrZ
w1nUF1cQ11kA354aFScPFCuK+i5PPz52cBEh1eiVLUQoJRkkA76VuMEeyl6OzUUUBND7EZ5sPXtZ
2JBkizIQC5Re78IUmqOTOW0MuidOIPv6+CTOEqUhsiirQ254mdTNvZZV4tyscqCKX3LF8vitTqu4
Yh1zRyAcn8xHTLyz7YkHmnXrgzeUkM3RxYtA0xaxhWP2BSLCDzEpiNYAW78G1nhkKdVCbLz+EIes
HeOVNNrZ1Iol5M0VQRLM+P411qFzDQvcMhg/ABq57cKAcHXZmUJCEeGG1c8jmdlx4X29t61PUamx
eT866trBBInGp4zJXUxclgRt4B7MhBHxV+mq5Cs11xtpWJrtnTDUUlKs0mDDJlnXQoS4tNMhxpim
Gm2Md8WiCSuPjrMdAD5NTKD1N4RavEJN5IMEkaH40FDG6ZZo8yzpu/a40jzmfOujnnVQHnF8u6Da
0HmjJZqOECUjQ5+F9VspTaE5+ZZu1WLbeQG5DPEJpJwGLyiuUEQt2/vBprTg6iwEenZvA3i7G46c
rC5qCFWjp4V9xR26EjgWxjeq2clX1hJauN0F39Xs8Bwxnf1Do0XUVQow8CBJoDCs68ezTY2U/eZD
ovlgLJ1Lm6+KyYXY5lL+eOwbYrPhRY85+tCLgCGQKrYi9iKFzqIRZv9WMqITmZl3St3oWklXxFoF
eE3FxwZWWdzHo+fUMU4jotSRDZJo8ABac48ju91QkQvkf+6XpGrg+clzG33Lp6VzzJoLkLYdMruQ
K7/3s0Z+ZcTpXbBcJIcMoJRrnzRKVDVBvcWB0/aKh9izG8n+PtCfrJa5bKuavnM8eyDJtsLvp5UM
6765ygXrAPOTap2LqS7zthIU30i38kcTKxISsNYEMozsSZ8rfTATVTPncIsMLR8h62WIH48xeNtJ
RHZN5zjLkzbVs/ah0uy0Y7ei6zDnrd8m951Jh0CD8OTleYhUa0tx0Qu96xV5dKb88BPKW2cd6J+l
5kmtW3SXQKI+1vueFUgtJ3fwgLXSO0odelNPMWrpjl8V88aO3aV7zhsbXqPo9YFaxadXjL5nsgNj
A1ZbWQd+jn4FdxkivuIZByEA3SFIAqmcyDH5jQ4aCK7rA9/XYhixU01Jt+ibpF37mhdvGA/RMB9z
MvcxjGdxJ9Az77Z2pvc6F8z7gHSQKNDt5mBH0MOJA6L+LQKSOnG80lzNVdf3MDtugK0kBBb5RdpV
7JwqjHvu6x/ziQOOcbpUusqoaavmTpi+MAczsjioJqlOZ8TDuPtoGL0VD5EpCBZ8xqWh6QNRmG33
X0F0RoD3NLknuCDuyKh2FVBnODS+8RP+/a+5OrlmFV5yiMhRWM6Tso9OjkIWKzXXPFpUPI5FF9dX
cpZ0iXSExLfL84zKjK2ljS+3i+BZdaA3N0Ibetw0jGGoOF714mljHGhDfnLqs8hsX6mpkPOZidAZ
2YFEtbM1yQsd5/JITmO5pTS9EAo2Ur8JshBtTtgjDCfr8Ehy7jwtXWuIbdqTxTB6U8X+g8ctkJxq
C8f7MsnsABdb8GPCJasDEWRLOAIdDw2NPH0ldPKxNZ5XOUM96wI09AKnGHfZ59rIb5NAUS+0KyKg
IlzObzlGx1Hl1VGqjn4EFvug7cxtzOkAxwh7GQuAlCjyx/CxGGXtSstnHTNX6A1aaeMzP2I+UtUm
JUXDdC6alOn0DcdiPdrEEeGH+M8EVwqkHwTajvUNuzSfDilFt3DwSAWo8NKs1wBvptqQdFY3mjwm
ugTgnxjroyYBzAs+m+N3Qnv5v/fEqICM1rQ5eYV2Mr4jRZwmxckxt/wfG7FzKs0+FCVpgj/pg/65
nMPTIM59uEvkqM4UEoa0KSm6BJLDMck52rwzeYL3LAmV2QDMaftN7g0Umrk6w3o5IVjXXr9BW3hD
XIWmpFBUtPhX4w58qUr3uDNcV3bvtxntdarf4ZXpGlfZaSsDT3gWQ4aNAT9rhbxt4n12Kn9YHJb7
+KKM5pniaEY8sPyHyQhTSTUyrRrGR+4mkj0ZIbbuJsRLTKnorl0gacoLAUzUPNgI3zkJ5/8X9Tb0
jmElb7YmBVorHFIM6BbZoWLN/XhJzRi7lNDYw7XrhUVDFs1tIIBoKDO9IP2Fh4Of8uk5rV1VMjTN
7QzSd8At3SikIHo85v+OoBRPAiUCVqARlf6HLWMiujz5F5ASFG5Wsg3F4J/3DSejV2gZ0dG64zPr
cLqe5sK8iOXzh8vkdMuqkNCVMrDQsmNY27eHvWqSd9im6wI2tsTytfNC9EzZC8qGZaanRG8hAVCY
mto/E3DMDQRuFhYcbftNs4j+1NVsRjBXqoGi+m4L270ujpwNdJsBCk2gXDEhhKkeuzkfYQes9ywi
JYpDsEIQikaHEkav/AQl0lyuKtjd30SPWJxn/T8h/oD/9JZrTV0b+ktCi3IZpxpC3Zp2K8Xrsqlx
NDFj4VAgh4yd7JZ2MB+8i77kdjwVtZLVKULzxNequQv3hosMwavpF/cpq6qtq0itQE3lWYoKTWqm
63cLs30n0crqYq2OtWN3nLMR76Xp9WHgq8294UW8fZh0y/BMMcymkDjXxr5FmnoC4eo9UrBmC7ch
ND1G0SZDnK41D+tqA0KKUt11t8eBT8EjnCexPdmQtwTcfYZ3e6PSue8tUy09URg+yWYTW4I7w7MY
ByldyJTjqTyfTyDtWKExp4qbXJQj30DELO4Qz7cF8qJalEZt4ydu2tXnod4lBj+tES2qpTr2D7lF
UZLNO+vsEYHq2AOEqzTdaAkl430SeWTDeFqdY5D2m/Y1LjihbJLJf7HD9pNcSBLlhnUx+ASaJFN3
s+6y5G08/cs/i4x6xhlEuwEM2Qp0pQ+OMM2Gm7fUv4gYdtreWmQ+Xo9MyuNo/NX1ZMgxHVQcX84B
MKZ1XXAPqw78cpgj1rXfV+ChFTD82bbPd/eihY5a2qmX/l3vSeboayj+kppLJxHK/9bIZlJS43DD
vsjrI7E9poOXPeJ7f5ewpOy6R+y46IkBynDQ2Ot/DrUwWr/xMPsqmG1NZYvJVxbcDEZMOxwCxYMF
p5YUrZg/Nr6+LXRj8Yvk4/My7oJzF1hR1rkLt6ObVJQVuUUdXvzSTKpZoSWRgPjoLI/fzI//SbmQ
efYEyNA+5u0Y6YZ8YdDn1bQA8trGVM3gni2ZsLvuurrVAroqDv0OfC6+0eeRvg1ENHphGZiT+uWf
KQDzRd8nCDy6RLRW2GCAu6TE+rRzMIvFIIjPQrfrsv5A0mYntGcqddQYyyJ+nmkuTyCcWswHD2le
36qHgzinwSPqpunGX0cWbNcX9YBZ+ZBuhcrWBaZCmLeGHq7Ntcbx8fjCla0H78PxKD1O88G1/0cn
kOIAEtittXf0sAdVFB3ISzT8m2JwA6VrW/dq0ylH/MOJw4lIIaDgPN5vzXJku5kSbgumxdVemmRY
CAGcYxB6a7pTYCO+KqkmrTL3USeQgHowKZXjw5IDYCWW5K0cLX1OL1OcjCutxxpAss5i++7Xcy26
y8z4gn7K5iwCH9sO9+co2VrOK34WpGVIdk7g4NWfwO5MLm5iX1YlMvGrRADFAJXQ+pXq4ze05l+g
4xq0sjynf6cEUesBhxI3SZGF5SxRaAyKrJFuN86E6nUHrEO0HHEBOpKZxqOmdquB3yX6YuDU636X
jgWlMpQcpXWHSyog4JVUZHG2LX0rnIa9PuMBQRum/9O7zWSUFjugWny8+aq/CxMh4zod6PSOAHhK
6yyqQ7ON2j4UTTNWabWVZ7ihUy6m+QOh0OjSqdodwHePkVyzjrzPprH8RXPiyT0WCU/saQt6zNNh
Ms+ZOywG+yFNPi/kPCq6EMEcHSMJEIPAN6U8zrDA1SO0KyjpJTAulht9INxFn6o7QE73a1IbOXTH
xFhx3moncE3JBWKXkR2+6oqVLi0b5Z5lQXej3kba20rdCp2NnsysMWehPwbc2ahzQb/6QRdeEv14
1i64zXNzg/hZv3z8WSH+cpNTcMO3ZqW1hW3lxMRFOWvb6iM8nqb0h1a4IayHzKjA3xaWQA7WtXJl
iQGrE17s6xhFLxsX3iRhXZbqX9T7/eyOFByhqeA1cRGV4SqKqULODgcUnXD3kJq4HMwGXqoAO7+4
fWtXVlwUBptBkKA7ivq3CMv4FGWnQ7ACckp+sOcpJlhuf4l0GkS851Yhc6eedVzt5i6f8FVg2w+J
EtGifSooQVEP3k7EdoDH7Y10ezNAza5Wwn1hXC4YBRcNN01mYSjbGfxoXEVr77W92d+xZ31ZtTy5
vGhVsXhURFrl5+aFJotaQ1zyvz42LY1N9dWR2L+OQrVEXf8dBs+UHCtAKiltfiTC0UpOD/ROfEIl
tHrFxLLuJ9CcpW1PIfEv0mGMhMMvpuF8WfxZ/4ocXdCG8KBqSRe+x8mLPNO/4gEbSehRjS0vr5xG
/sMF7ClbGtJmy1pGUw2CXfZAnY9d2zf/4OSAcO8v05htwRSV3oXI6Rn5hI3d10nJLtGzMIU44qu7
NP0uGGHdN2FCcIUHAbfoYAoZZBOHFUH/gizNCfRX07+BXo0adstTJKAkgjsL02DsSFAGGyJs5Eqm
9lzASypkGbIX/tIG67tEQxs34aa47M7l+NYPt+6BW0CkBYJ40vDvnuGH2LcMkYMRy4nvi8rB3c0E
7eb+GobQnpJQTeyyvlfNbF94PAdsuQvpHbvwf6dz7CBxREA6BA0iDKWAcMJ2WZMnGCa5tysY5O04
a/0MTFpP0JOhFke4ih59XBCrJhnzcEC55FMzfNd+3Ve8rW2TXmHHv+aZzrxwO9f7Q9CHHklub//A
raOsokaCBxaBmJRQO4LFSkNfzQL+VpHob+DD3PSVQwR2tKe3N631+BaGEWyw5GdV2BJJ+71UHmR2
X3c/VIZYvXQQYvsQHIhBdD/rLQ/MYMQMKrIq1WpaNeSAMuby4qHNuNsePl6cHb1QqetKZ8twFWUW
a2rf4dojARtC48lZ2WN5lda/P5YDZKiWwvppK3kXUuYH7FKOzkyvTAL1qQJ9wNFFlpduV5qxLGhz
pbd36t/ccVWXr3u0O5hu59rocqcs8QcinGLWOi2SWyocZkjbQrnZa8SbaSyHO4g/lz45oCYsvXtr
qMwWCOI0zHiOREjidVGDF3GAD6hX3uZH6mb1kXzkG28jkyotxTe7B7FtwgbY5v8sdYGhrlLNdzsE
UeV5AS933hws9RDY21p2Id1veBz0hxv6cA5/oGX56L7rZ4WnEkgaHYHpr/yWmnq10f6wbmzp4Jeh
sxdoXgoD8BI1CshDRmDPgV6oZhmibdXEhs9256P0YsB4Kea+C93adj5D94w75SR+mGpPqRFIPyZC
Ja6BzUIeLPC0aIl1nKX6slzlV/Kxt54fzHcnUjFdjlbY0cuZQX8ZPvBhFcpOwXbJsC/hgfziLeDm
DBFg3SaCYmDgeOk1HCCCbKo8yA4MuJft22P4rKLjCSiX+wirtPLClItZ3zp2Z6RthFujLsfj1QCZ
c9L3OSfwxVuSvsN8QGO2xZgjkNS/JWWICs0HAZxmEdELTHyoTZ4mGfy8N0Aqr8UHcYiyyMAzF6P2
2S9avflSUZDbUh7jq5ZnYKNea/L+oYlqh67qj9KzBe42l5B7Afvd1x18ZWqh+I8fdHnVBG3INPeL
hBzVmQfyUZlhTbtY6aNaIdsoxca7A8vysrE7eudn+2NAnfyvAw7Cy8ZlKayLPIWs1j4CSoRxjN4+
ZPKaoytDORKfA/vOres3/Cw8Xxkw1GmSV3tDByDjAmnyec1PLZa3ufKx2zOlCQVth6FT4lSCN7+/
SWhLTwM0GYNYJO7/rdnUNGYOrv3HXixkYrQmse16/7XG3R4CP8v4tttPaAlEDnrZ34DqH3cWygf2
3mrwjKmigBHT70lsVj6ACbDz0nkuXa58m8LObPBavyV+/zQBnmtgEKJctfdUuK13ne5RxHwiYrrs
P71HXWdeEiOqyLa8DlxaMyeZVPznBuo9Euntqcca5iEr7qiWlQnrKETa8rq2XI3hgmc/9OlVNj9N
MtbRnPkULfme32jlw3EHThWDRrtxhLcHlF7SX51v4ZS9yp18pN7walBYSjBydgBOeAhAWmg/h+WD
FPBiW21SFLvPAsk6I2lV2BJ56uSnldCPgMkFdZlOpOj+5px1w5RWE/m1ybATU+30+HD3BzF5YRF0
O6eVUwpJZUPa4nET7jIOp3e6Z0euASeTaAqwXZ3QzTCoOBieMmU/p0WHuO1+uidI97JS7gqn1t/u
4rehheBtAWgOwX+gUx37xGJTBYTZgddNu8EqLRFxaAYEu/zN6WBMmCOpj0qQzsTGhw+ZAuwc3ngi
pKVambDBfBJ+JagZCEE6/3PwoAGi0OMpDIEy7AD7EUpHT1sZuLoWd5uVPOQxeVL+JcaUBDbtwp63
7NwDRPtZY2t1NFKwACTeHAJeOWiyGj2RiT0pD41qqgWzNMi6Tfo32WT/kVtSHWVyIWbwsCoESvbf
egj3aLvPohe9WdUyIGlOoES/bi/y6vCthVnbr1jhvQppp8SuTtYBLwlFaJePDdTuUdH7vIvkkyOO
Ld+kLL3+rAECgvQEB0fp5Y/0RwpVk5n/X4eLQt1lQagA/SEVvjGwo07WGF5kHPZyX3oBlCf8rZkH
Plp2XLKMfnVYdBkPFeEZEbYVPTveaSSHF2Rb01GSkn+J3nV2PY60ggrfEd9Nqid7p4WqrN2qwT0O
AvCwzHJADZZqp8lpO8sLAiZPAEqbEvpVF0LFS4O7rY9DjE2McYdZU44EQ7LgxXCesovNJHwoyro3
n2qrKXe5pAIBu/+yZSLsqi+amLy1e/9uI6XUDaM2D4PhZ0eSJz1SCVNArc8DJK1IVskLuL+oT28u
Q1m9iJS7JkbQV/q6IV24mkoTsXYs/c9Tvg7nwkGz2IS30v4UeGAYp+oFQYllKfAi1eVghXkRNMZk
u5MUxR0ELXBR3IIj7uQfzZaIqpew1iLU4V3ZSwU1DXZ54+gpCu2w5NZ5bUyP8cwdGMGahKTXaPT8
b7HiMA4OvxNXpYhx1eL01P0KFsMcrcb1B27WwjHA7K937ORPeDaZywaXXMdJ/HXlMKmgAG1+Turr
4Bl0nHcreNdblzRU/Wpx6nMTjo62TzlCITvgAmRN+GXLLXCTsGMOCWWxHtW32mSiE8v6fFMaoPqR
Zh1w8qe4vQz8xiNyQL1ds10BUrotbq/BlLCC+FskMPwYrJQBj3VDnM+lQGeptmrvbly/1/I0NgUY
MrLvKM2oWWhioINuXWmwBgZVdPHvMgt2D2tn6q+0R7oUOK2yuAiAlVPP5LKe87MwRlPjlheL7CJ6
871+YYYZQdLiUBKjn8wGVoIfB0FxD4SNOeHE4rpCcE/r6shVbf8Mca9LxF3SyJnisKURup74v1Sa
e6KmWJbA43sXCRxTJHtXzfE3loD34hKS1tULeFAO2lGguIgs62H3fcqj3ooOIAC3JOUKnz3qi8tI
dbawDwn2PsCJ2/h648YTPkWN14AlEiwfTMxb8PofsdRQyTzcjR+jygyzELour/hgSADetBAhe0uT
uYFvggxvkb0gIsQDfCFhHj3VrMJb5YXwSTdVjRPuJNyx+gHfcFt4m44r5dDkGuxBCs3lm9VO8y3v
6pwH77BbG6q/KKjsQJJ2jRZILOvv6HrCznXsUgI69+PSai1CUlUghmuRL66EjGoa2xjzw3PpEKwV
qwzuBG/rsFoc0/YmoBCaCNhKO+61GNWofeJaWdr8psDHVbfSLUhCsIm7HbPl+dAHIhs3skgCG0t9
ajtFNwL85fX5i9U8/TI5mvu/r9ljOICajE7wQyB49Q8Qvgq5W7T1yIMeXTeG7C/ak6Xk/cISro2g
3v9CjefAaE/oQeHr81CANsdZZ6//vgWBQio+jEnppFdqE1RgLG9KLXhU+QXp3tQ7JLZcxMfVB0Yq
07Xlthm9vg/AMb0bAdFhBoZSz87g4ty5kUs0enUjvzfTyN2jpUSsmlKZCOBayg+vEXKXJ1G/oj/D
D1LWcDfCFxLHLPZQYHR/VHtQB8ZhaCzlzb3WPwB0DX/9aewOU5tTlG380A7fPZqJ+HKZ9MTtgiXM
u7NJZp+nM8hnWu/MG/g1t4LSO/EFRyrHTeNZxEHvrRAB8r0iB+iMRW1zIeKdNBFJZpXF/IqRvFtf
zNQdWksZRrRXI9jzmO3j0Sqwz5gi3pQe66zDJJWznbZ/Z2Elpw5lbhtt/Fi5cVcu8iGwMBMMOIbR
hGKns8hUhSDwp2VI/+3Iznq2hxHrhrMYsvzNctwGFDY+DdSc8usDJaKjKCoEFaa701ndZa5dxEny
gyvN4nL6mvBisdXfRJOXXJ8j4Mwifq7/lmDrMd9eV8SFKdz40oLtoxx8iU72NwHsSw5IYJkkPkvI
LprvOT5RayJ99IUomD0ID0aY1/HfyW08KJGSKQpKh3ZAzeIro4hUbTtsyQ3gzOQe7sVsOL99KxKZ
3mh6PGyloc1roHV5aNO8MNhc5lgKEU3IgUErTgLyptRzHG54l/RTG539bHS04FgsfeQn2awph1oH
vgfAyz6p5XZQpYepiMhNdevDtehqubL+QPsfC52QdKqdRa/2d/Rr2PCJ5AfzCVW5jZ+V07R9jYbF
FLy594IiN05FKKDjRRoMzT7kIxg+RqQRI5ZQcQAlmQkL9si3W/lP7Ayl/y5UzXFMfFkJbp0GUeFz
FPhNMFNGT7hKta20t6AiEIE5tdVYyEm2TmjZGPomCpKEJNasw2n0vDVFUhZbO99zeXAbJp+JT8ax
BH4n3d7bquWW78mbkbzVT0wyqHLidSLHpBOCAPTHDF6S7R62sSOenBZJuOqkRchHWu9NLEY65+v3
NvX4Ks21jz+LKvDVBzKKT+Idi85ciaWeI4FUJpESoWFyAWYfwItYEDjNmHUfRwC+FhSYArE+nTwh
zj1HTeZwq26fHMzGpGHN5vGG6oAD7HTFwjy9U2wkmheUYpukWE8hLKGJo/rIhburMYtehPqEbGLI
nvp1W2apDCkzTjKqx1EwXbkpa6/vLJbkD1BFlRaizpH2dqQ5vb8ym0ve2sc99PgVp/TbELk5DLxy
qPPN6WcLrNVhXxaVw98x0AgFw9aWmjiZkuZ+JsGJ1GDmyjCj5zoLUeboWIEN0HG353gxvu8XpI78
N0Q5C90KHg/WVrDi772gD0/WgwRTlDaaNbDco3POROSp5XNLvUqIngDoH2hF59Km7tRNejPcNyCA
M2+qy57R2/xw82ROLXT4FLQb1NCMq9Wv9s8SP1rrC6RmWf/BeTPOQT3DQJlmR3ZjQIGNoGRY/Pdt
UU+ZPWQUpKocorgrcFKfxlB6R+R9a5fFzjKXGeFeeOU6FDI1BGSYTb82wy0nnRQbWUblYIBMDICy
ARK73EF9cH3LqRvMK6uUTUMFdWK8KVxCOPpr9D+gZVbo5BNS+54rp+lpGGe42/b99B06ovnumI8v
X2eVytdkzix/38ARoNURwApenAk4qK9CeRzIWtQ2bkSYH4OBR1fo4KoLLqcdwz82n19FiSUbO7S3
tKLCuMDoF1oA4jaQtxitawJyweqxkT2EdHX/Ux4/gtxTHZJjU0uMZwRJQZgs0B6H4+ULKpA2Quzy
EemFjiyHm3y9v09MEX9SLi4+ofu6wq2CxoT9ImSk7d+2lZTqwlaByOdSMf4ZrBVcUghRuaL9Cj4O
zjP4e95fdVzE7dA7q8oZGJQEuAFKDHWzHHwfTQfA/MgvY6itYTt60GjyGOfU6VCqEoAo9nXX7PJH
qxepDTNZbuBRCaKjjGxFEXNs/dnIojTC4JCygulHImY9mG9WRZIiT1tBb03UJj2buhOUOz500VYi
I9EwcHET+WFxS4wNlLyHsXCA5Bfvi4/CC1KyFL1y4a4Va0GL4hP1JV3YlQeVicF/8tzuhJR9/2yV
Gz3nmP/eETTm9NKTCA35kl2Up/z0qTf5COmjlyEsGPBtUmOtbkZ02WXgyALI6GYq3O1OotOU/yh0
4gS5cHOmAGitIrS4zLMsxMGmr/VrEThBd7PSj0osml3u/9TCFHuFM3P3xWFvGASRxt/tcG6t81++
ncw1j/pWJcK6s3qPrp7LKUAXF/dSihszt/ebKISMqbqk2Sve6Itv1Ji1vKXAtU1OKWr4px/tS6Hp
ReJiBZBRuwUFC6AT77NnS3W6n2CUZdI3xaoZxzuJrJ2oYu/+vQNwE28zbC+9c6LFgvr7t/6EBRPn
gkghKG1VioVUpVeRv6WjYfzP/ErEuVXOwtTSjkO9BJm9Bp5hfkNZnt2nIelHbSsi6d+V3jSUCiaC
lIK/up9fUDVkDRM3XYu5JBcMbcVN48+ryHJfwGTl7O/gG7dUtDwtgiyVyFvNtsLEtQfN+NrBjSHy
1NhTUez49l4CuPxP+eQ3fr/x04lvFPOUTjzDzrHA9cQMpoHhOaKx/QpvowklFEDmPZq6aMudLtkX
RopB+If65YZM9Kt7RjULfobBg0CYKBcX4fpq2LOv5czlli5XmB2fOB15JP50uFeQh0gxIHWwju29
t54M/w4agGf5K3cOz//7ShjjRK+vH0ROdJpcx1V+QukmtWQsXVniE/WUCH0a6TdtJBrX2BwuGoRz
OUrVhioGBJStD89DhfIZ6Va/qLuJbHwvnjUmD+ytcytvJSV/85+9LK/Ko9rPagitYDDTIDn0xF/J
vc/1otGlhCesSKh1chqG3nSoS55g+X8Gr9Lp1tyGn2fN+pWMRu3SmiAZnjMXmLwl9BQ4rSuv3Bn3
iwtuZGAsm87Muj1pizji+/LibCLdTsGGbH8/earmwDHbyNzAnUuCUvOvT0G64W7zfD0hVepMBg8P
r5ncykNRKqG8z+aK/ok0EhecOBWvsrbmv05xTln6kJ3kg+/gZb+j4sSiKaQt75/GkotbyjdBgI3v
m0tRT71t91zKcL8a163R/ZKBj2k06ANaKE5B5f6uLXawZkbw4F4rLAHv9y1ajfhs1GE0vg5pQ1El
WaqYPa2fE1aThEjxZu7/HsQuCCEh8izqO/h/2JZESE42mjNkk6Rggauh6lx+2l453m6PMHgskFbS
rwrGaHh+ZO5WLqLQjWdr0ox5zFGa2jwJa7/PhEVAn3bHfPcqH1M60zAzxdTt23u28HWEsf/yF2cb
Lob2mhSOzQ1+bKeXmd7URz+GEEXIR2Gjb4EtqGgEwLXosbyLR1R9alk9qTlTxFCuGX75OVOSJdTW
6J/aCGviMR7L5pQsFfKyeAZq1aKd7/pqE4AELLdcRKTjC7WtO5nC1wGymFujxwdRCrSd9KXufzlQ
e/6YUZfCtFiejdYSge94ekEMwtX1AddJ43j3xPzUGSD+awFIcYjozDLdUL9rG0soauvMiXDrwgRF
ax8292vuQ2Af8QNUQM/WX6moFFiZgI4wmPKBTkXplktL5S2YPdJZCFWiTImbgPrEUcCjR22Q6Fqw
e+ZBktki5LuTsaqxvjNIa93Rc3aQuMqHt2Xw1sorH0BuV+zH5BWCHhZV5brIzt1Nbnzy0qwmOS6x
hgYr9RrS+5FwirBBon41zZJqC1mMuaq9Mu49E0fGZCEMqE+oMsVEta++Bu5Tnqjdblp/Eoe5zb5u
yt0I3z7sk6/6kn1E4oguEhwfnA2nJKhk/2Q5jGRlc8V+YmY6gCesTyEBQML5RRvrnY7VaUw/Yo2A
LkIzL/cVVBvjkfWBziVA/Sq/u9dIpJLiTuELu6jyDq5Sc5vfi7YBFVKaHEL6BgWGFNsdg7YbYSR1
rOAAPp4yC62ydkg+AJnkdQqxY45MsOCjvC/dGkdOffqcAk0ghEmDXWUGMXLhEd6XbGLX3v1K7zAd
cY2ygNSfbGi8JvM/DZxmsJEALdCtiQJiB8RXQOl59QlZZ1gCX3xdvrdPMg/A1phE4T4D8Eg3xiG4
YPcKRmiXu8CF6zf8X9fSn7SC7m+5HQQ+7y1kjn9HNxJnwbizv77V/3baNgb9ZfPe3gt3Y/eTqs6w
eb1R59I/PseUbQWi3xuqQ42EDr7Q6MBnBA8hElzd/2LZSQKr3cOvmYx3Rh0UjQ5CiOU6RYbLxA2t
NZmdhUx0qN8oqQldd1ctCRQrz+sTOWzT1HVCXE8OuDLdXXu1hjkXMwVQtCTwmtcmPwO/Zc3R1SMp
/GT2KMh8GGZDko79Z5TTrmv3u3zm68nkTadwyhYI30Qg0JwlOndFn5wjIW6rhe16Dob4fZzPr40E
KEyPDM4hXqn4J2dFommO3nCiAMcSptjTpeBc/Omdm9GJfuMqyzoEX4sT63UDC2yRLbYBAuy7SKbm
VpIQovVYkeupcM3LjNQgF7+YJbRxUCOSC60S3VNuiOGuU1AMpeU4SDGbsfCQHlj/IKSw6cziOkvk
8DI2zqDB4msCP+Ac4kS4FU5QbbJbyotSaYcEmp+Dwwb/F+nm0LPH/mS2VAw1Cpxxi7evRNs+zbzj
SY+JhHXha5L2qwPrNxAS+X2qGFATyHQ8LLxAc0SQMyd0eMnk+uCHkH03A9iFGIJ63dBbdSi1TAu7
JayVwASbuE+bdAnRnpjEH9yw2+VGZHhKE1ji/vWtHNoV1gg1CMIWmm6uSdccoVJ3Hb/D7yip3zFG
lJOWQKl/0d6+jsr/HsQbpQWfgQezydSsUfzoC1S+1h6TKuhtDCT2MmYEhGha4lnFv6nEYslHjDlZ
TpbBP9720UXF9kQV76ZByWGc/+nGfqb2eovyBi2U0i0kdZ1Z/EGKghjwwDbwDw1/vl0yXOdH+yMl
wyPbGCi/gt24g6YKk3jbSswZtw4+ar3UbdwgH/n/VVkO3bXZoE+mRqOWbDDxoshSiVGhbz0AmWzd
iSONuFm2EY7ovljisXV1rWw1hjS+8Ls8q5dg6ORuPuRI6U9lZ5L93ZjxLkj0V9gfdJ6pz/UMgoXf
Qzd53GMbK9zSy1sH6wmJmm4U2wxN6XKfF8f66Wi4JF7bZ96BbmrOnt6vchUwX7aHoSkS8H3BBSvr
bVOaOAR2LSyE9ezbpVQTJSfWRGNbbGj82Q9GhdqY2QrwjJMMZB415wMLukJ88+/hIk3lvwn0nA9z
jNmmiobvuC6UKQTt9C5IZvObC6xc/BZ6Re1hekKzICqpYmq+jhouTPcKhCjElVS0OjEOG2kYDL/F
QIumTaUhT9KvZeatxK0oWqhUvhq6S9r7Fx/qw+ceM9Nix/B/fjEfqUDd1GxHaadI8CH/awxtbHfG
Agx5mbtZt5HBKWNkKr6bw2+zDDtIH0sIRBbn9ZA8T9sT07d4LMie7OoleFmj87PzeSTsAv4HyHki
j6Kd1CQWhwi3qT0l+IIOwqqrXYwnmL43gCt9iLOD0GlilhsNBAHbk0XwNQ4Qd1w/muMfkxJ/QlxV
JHFMkH3cX5LzwzukduNIkfjwpcl/wKgRMmzt+8sBwqY/bW4ZARgJCuJpL6lwfQo3mQL8ab0qZG/j
kN0WJiZXQhg/c5vMHvLt8cEX2HLOgFHWarxaMJ9RdtfecbPwIPYfDW8b9VNdCOfBJtsXMIOc5o0T
tmf7lOC+QTuescP+Z6M3LWGqa7v8pGYE8WamgxLrLhPQ4xXogyyRHTiLWn+Ia0BuE0gwnl2jlAwq
D+6xtLqOnrHizwAr3TZ4n+XYLwayejXViC5BV7SWn2ov4GLv4F7rBekdiz1E7AjHfRwHLU/2YBmF
imaHKPKB9xypoIaUqmuSTHWTquMZNwmzmQEp3w2lyKLmyR4gOVs46PDQ9dxTeb6URPgdqfM+78Ge
Bnl4fKpPPVlSI7k2uyRruKpLVr+QB394kVDe/7u7A5EmKBihOPdmGLAGTwXE5CjHDazuysUcM7Su
AQSWrUau/KCCZGUJEqxw2wrpTCZbI1S+l5nwPHitjy+5pzhEHp6DRjlRCTqg4PBnDGyPqnwjRS3L
W3rYOM9MWcqYFz6PPRO9qC6toozuRlbinjqwYKo92ankhcFbdsQ6hpNrIfp3KAWULQvYWGXYPcNQ
yqMsHlIFhAuX5BnyOZjlO3N8iMNocIzzn+OGlMc6XNL8fgT/zkVkQcUYYZJEpiWNTnDhyjaz8gAs
VR0wn5aLuowHnTl4phFUC3vRTPGh9DLVvasao/nhlFF9+4gG3B5g+iTqMAzb8hPoy0al+rmK/HxR
kGOfYjTl5alDV52mr2S/xhbHZHfEYB75wMPUUb483zS06BFto07BLnEaAl1v/sVae2ptYjZWQ/eR
JpPgSEjpC86OzGHdcH4r3LjK1IbUTu3PjIxSE77NN3/qZdpMvtkzsP9YwHOuTjdHeaKU/iESzyfs
2ZOLvUJGTEuydSpNfa05z00Y4YoFZum9iOWQYTqNrA5hTdsW4uwajHOsO7Uu21hi2eLHCTo5HkKV
kodVzXbOCXOJ3EXl+hZFEN6EoFblL2Ej+J0woVB0oiJM6MmQ8dQ0TsqF4N6kptItJ7xvCdskRNaP
4s9dJpsp/0OYgwsC3pNhr/eaRBovLUGS9n/P9w0RBMkejcmjtT2s3OVg+kVdWKbCTI5Lq4uLJWvc
CyB+jM5Jer4Ns8XHxfgktGdIz7fUP884GDXKkTV8tTJeixovIw0PQDx6eyGtlwsuZltuf6LaPNJH
kSCEjgw44CnKuGqM/lcEugyNouY5PD8iX5gIvwfgCW8xZQOydcqkllPGs1cRvmHPjmGB9xkX4e84
r5FPbAQD3s7p8foQz2M50/Aq2lb5BHsiI0N4BASiPdoJYiIJG1+Lt0JVuth3f7hjhTKb38VhZtNa
VyT5l7lpDOw1M3KiGhm6E5pdRrtgGWVY/YpxAmSKs8Us2Sc1E5k7JchXSnP2jn+iaY5lwvIBrNTR
vBgJWM8HEsGbJUpMScNBDi3a1fK5AJX9IZSbnxv16V9ooqgf/o+1tav3p8QZLMA1i4fmN3xBgT5i
o5IZ7f3YIJ8zcembJxG8yJ4UEIJbj3Q0c7pkMrP2n6463Y0/NMWdMSEVdoCzuDkFT2DyFiwUlJ13
jgp+2o3/R2Qn9hck4MXSBOl35VtMHu46ENwz939P6wI9oO5kJEZ+GlF6j6OUsqARpa5mpkWHZrQw
LwHn6mWWYH6pSsY5znseWnf8Z/vxzOASULPWiE8WiosDjPu1DtwLAJrgPWliC3c3PduS9UBC37mv
LYVF8n7WM0dPKqR4uGLWBn5phBmGSAeBn81r825uSgK9jmLUG+X8cffRIqJuScbMHzO8VmtMJal4
dXD3wwodLUHpxKAtsPxN8thNnR2Uyt6m8E1/7XuKMbBZgWsfMptDBdY5XxbE0pE5MUALjrv7Z2ML
LRmnSpeovLHdfoKHOC7evJJ/maKAU+2g2C/77poivXWlXf2iJkXCAuhqpfwthzg5ylQH9qK58vLh
RXFZJitS4EFE5DTHR9XkTnohqIQcb5esI/b3xXgxEO/e8+t+WNkYQeEpn8eqfk8wvn3KUqGpEy4u
y4J9Yux4eIM5lj3rXNddVp5cpmrOW5xzkBFMfFVdFsqubLOFCKGcPcWQQWQ3goWZYeY0wcPRcv9g
UoCAm81Vi6W/EUhaSxm2VUlwbldKYpZw3pLZ2O91gAft/eANm0USVsq9JAK1cXYYnhdYm6zu1RVC
VYBditHXnB51dshbxHvs0ZmdyyvHtlc+gIVma3WHSsbst5+S/iifAW0s50LrEs+V1Qh9Pc1fUHnA
0u9V/miQ3VwGr9sSkpixxZ0QBJwWzVPAsFZpf/+7v1eXM5SCG2UqkvJihW/VoNbWu9q3OHNfewgU
eS6nn0YokhL+9tuIHUZ3cVKbTcc1t1qYz1JvcDePr88+mwG02jkQHrOeVm55RJAqAZLuPwRqf94W
oTPST8VWDWMxrUhHjgP2xz5kzGEs+weQf1vis4y2ydFTPAMCtRbvDj5IjOT+cqPyz7ENeWLqy2LU
I6ANBW60YnQaykg2t2rw4cLnzFYua8RmFq/5FqP31WPyPppJ4eDhdw0kDVqgco9tb3/i/cwq2O+B
lUmI0OhNr620jL3RoTiBnIv43Amprrl7XzCXfYpK5xV4MDoimo2KkerX+yfLDKs8BWFkulZvTRxe
zuJylP/sPChkd8yxnBEfyVkCFdDrfGzqXY5p6U8/kLaz+yknMuUa92Uw1uiHdPh2JGbCQwSJ8mHp
xYAULgK9LSovtuq9p2Pcdt85Xm+Z4TN4/G5eROVA16v+uFMKXeljxZv4ObhmmOF32hFg8ltxRiTq
hT9FMcbQXXrsgAlJqAPdwLixjymNp+LR99QGeRdcUeHQzkXk55NETVkt/NSs2APE6QkGVygi0Qkm
2xPOtJy6Nd3rSodhSCDG8OMVPYdJ+QMfIbluoANK6sxKo46vjn6XjHYLlTZZZIdfYihuwfsZLGbz
kv3f7i+DeEIJpGdHstC360BTF5U2dQaMkO/BSTi8EdqbpzmqRfwyks2xfEt3WDYhINpAMDkb63KJ
LfzIPZ7FdP8/4QacKkUdIE+DJ5s4+MGEpfUsuq5iX0B3TGjXtloGlmc3RymypiTI8dxL3C5UHntv
88UO3Dl9+K/CbobK/BPZPIjbOwqXqMDvagQBIZJ7+qVRhMmg1lQXYkXrLfV6gOQIXp2xmbhMR3Ey
6MbEBxtmdRhhen04VJfPmIfS7lJeHRwtndlsHtvX6o0BfSvRNJVdHwO4IftSiCYlDVVqTI1ZGMrM
+EEU4LbJf6Zqk2edK0CV2ISRFiEVSOvtgb1N4wwgROW0qU6dceNaboCSYe2bhawNUgurxCXVkQ/J
v2wsDbicz3KIubv2PgJahzLWAMn5P4OfcooLW9+T6mcd0hAWB4iuehESwo7hXBAxXm0OUf2Q8WIL
MxhfBOIzRz+6R0Y4BGSUnSv3bTXl5EpshisgO5UrW9jriJ/ClkQCoTzBeGNwfx89SDRGZFDaKo2F
kw3gum5xLaErgDGjNWUaGY5tfIHzcaWOYdqFNl+F4ssusReaNFstAOia3d81BoQNkXud2ZijSx1s
TUSD+2L3I7ULzNrhlpBN5zvdJeDnJFYZypFvASnoJ8leypUWJ2DTgeHojVdwKWDpzlXTS/ZxL49a
cyvp9WflJA1Kspn/kYT3YwU+Ltl1150UklS0bM7/uWrCO7nYvsut/apk+mygyb/GpEpRDaKk8aK+
r1REKIcMyYFnkIjaPSWur91D2gIN8BEK7VqMI3W5qrx/oD1rn67yni1koOyWInxG5U79z2g6SCxs
8ou7FFBhCEk8DBehfMnSGcJTc9z+0M2MbjmrjdSMxwUHKyX7n+owOSSH4g4m4pa8MaGCzCoiB3xG
XZehpcjNozO2fsMAkh3RmBWtA2Cn4B5s3XsabKIarW4xv2/NeOvk/CDQWP6miEUer9M7laJJ1nBs
b0vjpXKQuzcWE+x8aBbaaNbaCo0L3ofn/RfHwDqQB8NrS3fhDW66I9XuHhm2YOrkcK2X1mOdL5+J
Sz2fAMIYzSxS/054a+lAd6CozFTkkKNIvgBDNk6KZ2jTq4W64FsZBCuumvv64qMZ6XUuXeeyafRX
K58PYV6vmIRo2g44ElAGgnXgPo0hMsJheSV90WUI6FF9DBJLhehrTsD75JVKe37VASIlve/FzRv1
0KLZgbtUI6jfH5kTvQ0Tfla+RSkkZEozwVrHurYiwgOkdC4mm3ALJzXzUacck+6ZDem+vOM42sKW
rolDLhFPp7HzDTcS9LjBVzzhDF1J48NGdwzRXgdI51n4CRChFiuMsYxx579g0PI909c2mGgBnbxx
niaC01imJOYP8fgx+0LQmohtFDkiCAS4pS/nrj03iwZ9pKLuMkiubWKGXfxEguggJRIvD00Vg9gz
3NeaUZGrTuMFMa/A12LQ1oUiyUxjKnCT/duiZugfwFzwb4SVGqehw2on5udjERajEomJ1XjkpMi4
bxEJmzKuWJ4MAwnwd2mZiZFhoACKBCm4ILrKOlMbEL9M3Nx3wJ52/OkvQzeYDwKw+qDiLR4VoXiS
r7IFy1/n/mbaqLLu4L0lkukGqC0KyFNc0K872Kj4BIJuLKKHNI3vNmRYiwLxTmmlO5UTWA1PQdFz
MOaVcokKj/CwKXB53LBh7cNDmsTpchIUmW+RBergCiiSy0cZv2hXr581682CjsaFoSoOKztBPW+U
rZkrQnS8X6XUu+u8ILyXKhCFAZybDbAjxS9J2xi9i4lwYQ4tBFWx/EivjRzA5rAHjJI/qAzbfxsY
3Vg71+/sVmT0GiCXTfXQFZSFX0l3fqfTvVd+h4N3MMmLiIpjAPxXMQHqx418j2VrhlkHTnsboxsV
2YG0WKNeBqTSF85sVtMFTmp1GzNODAk37AU68/Ic+S5ZpTPAim71QxWzEszPThJz02jpdXSZkgdn
XfP4Hns4K74euGT3l9XSSX/wVJm5xPfzCUBUDOleASe10MbRD70riCgUkMs5PwGXGiEUxkSXnSBF
G5cEq4LInNwtAr9btl1Ebm9WhiINcDyuCerCTwvbwn782Ww4WmN3Dcr0rOW0ALjDVOpBq5LIFidp
b1rvFh0BAk/9jTS1DxsExnrcqp8pvGTT2dbPz36iYK1L2dclQ+e76w3gwOmQPPNLWpSHaB8Ias4R
95DBmthmTK9ze4U6dA8VUEvsdq8Dk7/VmXZvQtk1tuQpgtoePpgbP+w76ch9wBXQBTmIj6V2lFwa
myD0ExWcAp+VZ5QzOHR4AlLifi2myzRyUPlBXmxWpbXS+8+qrNb2RRn7XbSV2QBGMNwd0So/6I3a
Ec5N+qiNQashoKVHqTINnXoEeEa0V798840fXt1a4w+XcrfUPC03ykVZbENV3/MpTLyvNMFeiMd+
ucJghEo74cOjZD+QvdMTTSh1iKjZ4OSgDWfV4Hz5u3gT2XqwD7+qGjl1XU0KbPm1w2tamJY+gEqA
KifQaCNxpwiZ9cLYb+yHJOUaTHZ9Wxm6t3I+j2XTesQjIFwuP6ORDaoG5PIgtiuyAQ4WJshXTZ7E
URgTU7vUuKwYvHDzeLtO2TBidLtX1GFPUcs1BNpSIKSnXN8t3RyxzWK5qJFKtae/47rcy1nCkYEn
OiUuAymcDBOkVlLLrWCb5aIK8FBJ5mn+JIyEAk8zazujxvJzq9dye0eNLkw9OASwxZwVWzMbnKhD
lKKQ8Hx+olSYFSgTB+7xXgLWUG+DZ2X9255yfS/cmBok0DwTAQBnVsEhRhzb5oZ6JmX6AiA+qpXN
JqKOIvaABXgrXKUMvrs1YfoltU+5L8YRJzg4vf/JmmsaYGqMSq3TKy0BpBoDSLSCBZIAxwE/1igo
WGSzK4wAWri+GY4N8PyX4mFbDbWZMPRel5L+7oSs1x5F5WWTmrQh6iejD5+Wukp8pIQX6SltN8og
YA8zlCNuutH3+wmsIKCTLsv6JxF5g/KZjaduV31WmHvKiaLz4Ode2A0nPIOvd6P+hkSGAAbQJV94
mPwmb4XlRhsaIeBIJqWYgVNdxGoabybKGzYwZMnYL+JMmYz8teQz7DPxbz7LQVSi1eC4Q99WmWxM
nskhoEz1Bq0EcJoJccSiIcbVw2hi/K5uT/Szpg+gVlwv+B5pKEtNPZd7PPrBs6v6sGaEjYm4yvUk
iqq9E6H3uQ358MjFu4v4gDM64go2Bp2pmDZlzfPJ3PgsZAdEjt6lbbhqOaEJ2IGTPOYw4kvCOMaQ
dl5Dz4MQNVZfqVwzah5z5k2sp1Ztzp6EzoxJE48MZLEY8iaPDA7p0io9TOrf8f707qq14hwKmrmq
lqDP4lgt9zbsY4ljLGj+eY9dotMLxebKt+jfFHRLIok/qm0XgMofLv/HKo+wlW3LH/zVE3w9UcJQ
d8sqfmoJoreHYkHalqCVuKKWLVG46zKtdoEw3vneAT8Q2KR3PLWb8hRuL9bciYo/uL1j+X7a2PGv
GX/ICh2oJunTSMxfSA2kYrpLSnMMHRZBcJ5frWB2cq8JbP/lNypqT2Uj14WZpeAhDdpovTuf6gQj
b4N+uSNjEdI/Cd+fln6HdW+ZHtD7VeztP3mzTgj8fqlfjlp+N/BigdrZq6vfPTeYUyd6bV0ao18M
zDEittGvBhW2X2TXpRwoypvdUEtKTbmvDPhhR1qvsAYuQqpSwYka/zKZj+YjYktwodPsQG5SYdih
PVjQtUXEOq1aWGB2wPml01SXpwtm2MsjIdmVnE2Izyqzb7F8DhWR5OFid57Vkb+8Q+i0Sh00PWS8
AryUE42Fy+VoNsKBtpsZwUCntaRxGiPwZTIc02ell5cd6Lzku/8w4zs9Js6/zYEWn9lFYAB3bhee
Ms8GIPM4Ga8GQIXqC5iQBQtMvPVQ59BgXgGcaLTBoPa4E+IwJG+7Ew8bfTRdv8MMcPUbbNNA9ld0
bKyYWNJoibi/ukqIrWTc2Qaq866/5EfCn/TMnvtzY1iSfIloYgam7L9jIIBFtXueTYDkbECkRYMZ
p/oN1bGcNwXyehNEn+LV7x6ldzPqJ8YVcq31Vx8Ae35MLqp39oHiO6c9ZSDTXYlx6pPfBSBwFNxe
RPHxQV+a5O9sPUgdQk+Qlc2sXAejgr6AnHUMPygw3JiD9t95BHx1SRsy1AoPK+TelnKOrzlStX6a
H2Z2CtVwrs6gLMAxaJLgoMoPv1PEMU6MXYLFM6FDAHL55605xmNuLvRsx95Z9B5/UsWMrC6hTiQf
RxtCT9zPUym+EIpG2yajojJhRJ584LlxYL52/KeQu7wvfsmauV9ZSHUp/JYaT9mNyzCaXEAi1Gqz
iRTUvdon0ZRZBjXeY1/nOSwf1fDZt3+sGfmmTwAHcwlUko+r4Jj4KmcsOCyeVUS1vpR4mcWnpxVg
R6K1YF5VgCM6tvc8oRczLw9BBcQ8qGzKdCUdcYparFL46RpSd+EaAxHyMbPJ9s5ytYhbilpPh9Gg
z9Ys9ImL7uzxVHYo+WrSTcJxm2Nwtu61AsWw/aNyY0UiQNoyeHTrs5vEvR+D0igDN8VkPXxYThSt
E+SB96nMZ8WddmNMKV1of9PLDaA28GATMVqN1jJrFYi+3PqU2vhuZJhCAvYagW0S8C1hNtw4l/G0
D1xhhQSWalZtnaMuSaxbtQUZxy7AxF8+HlylEHBFYNZ23g5ojyrnkhxgRYNNACQ8wXP3RwuhVFWQ
ws2tUs86w/s9AZkOtVAwWZnqBhVv7Lbz/SJd0Ee/Fg7IoGZR52Ft5yaa5DOdUfkEvGqtPO6wtsUF
/jTmAqqcdxkys/qXwOckWsstcMzOm07k/7flFkyt2tceKc1YumLNtjUyzWPfzQrdZUUAPp8IYE8I
EsFzZzBWk2w69/Jhmt5E20CO1q6MlfhJFewWVMT/GdIMZaJ33IXaTpERdezf37GUWmyEN2fRoBdj
7GnIKrdl6ZJEZicjfO9q0ZKDAKjDVuC+4PLHtE9XF16KUQ4c06eEVZOvgLLLPuvSkOe+QkHyQKkH
0aSf69Z+5zbXGmHsCqjyxUrtGhJx6eIrgSgNsY5MSqkOBxiafW/+BPPKduesQXL+FkYUmCMohh9b
dT/h9WjBB+IXJzNcvRy58JaN7nLl0hI0q0Q1e+wx1/2uFTxzYVkQzSDUfW8U6uWorBC4zHUG8QSm
My6dk9To3Fxt3GOz++/Ykz0jtf++eNfMgS0k76WJKoCLkACPfCVp4sUc5xGcYeAYaTBMEpsMZhEk
seXuzQD2P6n/++4S+NSVeT0KcZLQcaoYv6AKwJrl/wgcIjztKURz2Y7kkVn7aFGb4rdswjwETCxM
BPiygvymmtsXGaWjSZhHvFekFtu1QTHvk/MnCy/3btB9ltyE9IuIuFLVGEjX4qdytsrxipkf6Kmj
3427/GmF6TDCACAdlLzNemTA3GPFau7YBi7y7dD2qEWUS0vZG0396c6xOswyrDpscAK16WvHmq6y
1fZQrkhFCaO2PcFaqQjinjQBUTQ51CaPBSylPcWjUOzBsjWwngMsKiP35Z3u2lLGMJKjF+GyDCop
y14Nc7OdP3zvvFN0LUTdMRQqZoWJ7LCRrTSQl4HOqnoKj/BEgim92+mcUPwD23OOkqFWkVpW7klY
ptJeoFRhW88GxefzfHuH72JbBkcyK/4ktqbGq4CxCYh8P+mpASC7PmkpH8/vOU9bzhujTd6wtWG6
2C0tgKtSPsu/8YSMphcObl8IS2dERQMWSP5C7F9LnWtTYkNEjFx5Bn7AgaB6j/v2oa2BSBWP+EwI
7VSGTltTDuS/x4ycyUlLNYidX2jN1DTkxbMDeu9vZqa6cKSKf+aJd3awMmWvh8EXszn+PpZynKnS
FT+zyHybvTbOUwZO31yYjJxhMS3JsQYggSCwwinfgy7pTiM3k3MqZweNtqNsqYzJpooFbMfp8bd6
Wq7tjAqXgPvWCnoWMEMuCZbTsA3AALSnaqYVNIfBcLzaYqccgz7Lq6S1QPFRcWn6VZAS/SeVZRM/
vYJ/D7k1n2yHdB37EnTsdDDw+NiZTBWOsCRTD085kaeb6vNSmf3W+jTWhi2XfRZajm4lAMD0OCa4
foZBLjYdUk4JbNgBRyA3epGNHphzYbDotwPcRzKrMCLdQewe0ahiqsT40B7N3/nO6T/5pW4cRNn/
5kyTLcP+3MfoedYnXegxrT3ArQS+23P31a535Y1VG++cnLC8V+Dixbv3yAqhCrLAXgFBzBs2747+
MVHMUn1k2HLKjkAiVjaRWcdDbSEC
`protect end_protected
