`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
k53ui2RDnpKDA9y8egf9N2jGP/uow3RIkh0jqBq9r0iiBbnjQjgmRl2a+3hurEaZKwpv8KsBSwcL
DRCxkws4sw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VpFcr01I0y2Y6jvuBmwnSpz9ElK8vRUTrdoIivebKHvHCWD0dikMvwHf052CGPLtfhI6z6XIpXlg
2VwJxfuIrLT/2vineeTdDuDnmPjaESfv2UN0IQ6vU4wc0h7yvIZgq7LPrN1Fb3cK93K0Sx4NdaSt
qm3j6+LSr9bm1gZfhLI=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nGmKOxFd2VNXuaI59kZTTUcb63fGY49/zSFap3Qr4JgxbqNMrIVjDBELW0GouW3N4gdu8GGZuIGl
wd8pTwAfMOR7TmOMJtD/K4EvKXTa4eEz0gSFKlT7SN06hm1DGKrY1YPwZ4yJD5XqKLMiLsiwH1S3
PQTaWrGEIt8HOpOZtyU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ERORbvuCv4xRLemEo+wDDt/B2r1U/1e28qhONHEdnrRgylQWbrpD6sZKGEdtWsuXZhwWBMvDcXJA
dPmJUhG+tEJC+fhPzae6/yiKN7R//LfZ9Jf+baSHP3cD6+0h4MaWvAdjgEZ+FOrtWAzOjfUh45Il
zzfBERZVdHh9L7vtREoKw8zVMlfl5kSlUa1KQrZ5zWfzUHaDgZMoPGZyM0cR4f4Mp+QWbvyWvSi1
r28iYm7OYC2c0M12o0RutcE29SfksWXPMbwU9Rb68sSEbBNcD9I2maivMqJnJwkC2nYRSwNuf4vd
2PdgQBQ8H41wdX3CRLktcdKY/6VltKB824kMOA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pCBtYYLNDndnoZyaOcYddtVo0fMk45yliSetWyoxvQj4Ra8SB535tZa3iqx5GnJxlC/D0p2hfvRL
O2Mz8oSxaznK8OLTEf1c2wUhuAIsPYPU1fZB2yuAVlvC7O/FAa9Vn7zByvJh0La5yNcxfRWVwik1
uPfetjZV9Kpb85fjV4MviCRnaNdWT7J5LSFBwYjtIOVHu4wAaGkV65gXz2+XpbrSMLuDXRlc41uM
eedPh7L+XLZmhvjsPs73cMawxYxMiZb9r3QAADWLf+p90vC6GyqR7L7R4LPD4P/DNSV5Fs+UheQI
dMZfO0UEjCy/I9vsuYpz9o7umkw+MC9J3MCnDQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KCW7MZAl4JDDMiiMj6VRXT1M+9ZJ4UEKA6BESdLZdC114SOFO+O8UjnnKpk2Fy2aAJQplaeJEANR
s0iuFFpA78FoHOF9e9DBI8T5i1JQ4bE8aYYLak8Okslr075gdCZhogcjh7fSYSqkk7uNRJ0++TVz
3Qrjj71a5YlwBnackHyvdi12TmISPhqpLzWyzkfPsmpmiK2GJejRqMmJRWH/1jIH1H/EAe/E6XaW
bjy2wYyW4dBgN1UmDdRpiqLa29BO3zR19VLleb2hE//NN32xriUJR/RKlIyUFVGSLwqoqWZNbCLX
i8S8MUj7C6Sx6DMQu6Mj9BE9V71D9rWE2aJung==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 648640)
`protect data_block
7luH2h1gAIHp+RUQV333acxdVbNnk+vZnYKuk6QNsr4Dx+l60q1L8wqVTsSYpiETXwsSO+SAGmqg
7kIPRjbr8oMWYN1rDlEJ5TgMnpZhp/JlYvdjMX3bpgpbu5iswF1s1uQvGOxOFW82VsOU4aMK+F/j
QrZCq3V4a+JdPUptxPrzYwJ4uX7EoSTQY4Mk5kKigWJ+uPly5EOQY+OiQsplgsszNaT7cKDppJHZ
fUvQWuVNrNXwuz5jMppHPVbbz9KlgeRTxuNsrvjDRRugsoLWXD5o1eaccXMUIRpMJgbcIjfZN+Pc
91F2RVYX12FgkihbVSt9GfC1Gfi6DpGEnahsyyqZb2Nm8/GpGh/LKabQP9v8qBRpiu0smkH8GPn0
i1U/eVdHa93GJG6348K1M6HeRJarAtuQxWqSXeYbRXMMWmQOZFo6suzlghR3z8RF2wnGUpaH0vzh
fASe2XiXRO7Lo3F+cZzwa3BFiwYy6Kp49tvKuMJaeVqQbZPkExn+pVOBTNpTLcUM0ALVpiWa4vtZ
nqZyUiX4R7usY0LgS0uholQxbYAati/qGsRz3WK1WcMKT6mLWnJkUT7Bda6ZGHxAS4b9U4kQ3z9b
UtDXxXVSKvCldtgZkNuTGYDIb+N+CFGw/qpBJhqlHGFcN/7jFJ7NXbTvLCIxfcFPUmNJgGMXNi5Z
K25iS3QkQlQIlq6wCVRFzCpbpwJKONy11mzA+4/d5GUYVuMu6pVTh+6G4zCRRV3QEIR5hmT1BXAc
dTOQcwnW1cAuANbWqOCRH08ewS5gEoVh4zaAXJUX5GAGMZ0eGUrsO2gbunXYjBbp11GTfMhhNQ0A
btk9hOYDoRUXnhPB8QCiwn+MJc6H1mv8lRyp0OQJ+E1P08o4s3LZigZb04ijtLVo+4ce0SMf9jHj
JDQVzRqfCrjv3zPoeQvg/j7+T9TzTshVtlSSAXaP7tpuSOTPhQCUTLy9PT0ACaPBahuL88y3H3ug
+6+MDUb4yuaNap3O+nN5tDUM48kZISUexshlVPCllxPMNXbCF45MHZ+qifxvKGN05118AIDBl/k6
91IX23I4HGh6El6L3GBbrBMeWsoJpejye9bVDeRA13VdyNEsFL1nhss3rD8KyUGPPoIfoH0kLOK9
ZXk5ILPlTZlfhPvosX3kpHSEK5n15ZiSXq30iTVz0TAgBboBqCA+K0639Ie1wnVU6uPFbxEOZdzV
yh05btQqd5ba6593Zo2FGgkb+bZGulsT6TUdY3LPdMIxRmKD9y5VZzd6pmm98FG/h7M1YvVSuYYg
mZUFjW/Jw79WUpH4w2dbB509PEX4Zr4m+vMJjgbIrENsNpQPc4jIUgiu/Qr1wq7Ey5hcy3SMV3E1
J/8r676qqQUirDq4Ib2cUZBlncjjmjCd69WLAF09vBVVO1w08Rj+RAdc9TQfwlEqdXvepThebgxZ
5XdVP7GbHdRvJpTY1yLrFb5bFl+hA+GhwTpNXH3UVjGfCBZhL9pieUL7U+vBnn2kPHpcn9gGd0Vw
sWIeEv9OnyTPuP+fIjOMnAPDnbZDd+C2k7WlV9YZGpb1+l23d9M4lJAEblWbAiVgcUHN47E8CBJ1
/wPFD0exN2t9kTSIQUSNeVhBnv5S5Q41vUr5sGocElf+Klx1z3iFy7mMyYcw8ACoWaT4lGECM7M2
HZwabIKWuBFNCVITN0c17F3+RJrF1CpgRU5oBnSIniTWJ4F52G9TmJcyBFgojNEND1x4M48PUQ76
rhytffcm1HDRRg/ySQ3YvoXzUKfQq5eDe6g72boiyUy/zfZW2xIn/e+Fj1ftYF5QZJUlPlrQOi7m
E9k0ZVIPfKm/LBde26YVI8UjmhO2DDrFxFuQ9TZxMp20wHNPbadK8B1Gz6xW0iJWVrn86FrsXz0/
4cG6uAltPQIyS2J20tHYgqAfSc2x72nYWIC2Z3L3a4UTO9cegnAEVs4+OstrKUEpiRyQf4/Xdxzf
cfzm7i3zQhuGCQ+IMDhaUfsrqhT/Yx5ySHZl9ILp9KMRlvJ5XIgYQ5xg05SCIBPO1jc41PDmKHTz
ainT2UMNoTR8B0x/xiDF7VX4pUj205MT1t5XkJQnzpj/WzGUOPbj3GET/QcJEKPgVvLywC8LOzCB
mXsViQFR5PeM9uRbPTGL19tz+G6xFdQgVUcQP0fRaQHQrBCJGd9GLFSdbKj+uSPaTHF9BzYSKjc6
0/5gJ6Mxe0exkopQFYGgSac+xCYbpVv//fiiOl7i0yGJBFh2QXmtEXMJSBTuX3s7IBG82Gre8x0m
/ZpT7jEaZpaomE8F0xnbThia+Rq/sZCAsWfCpMOF/e/6pTs4gFkRCKpCLvtxbXXL7x23/HDCDQ3N
+DYHfCeGM4pN626Qfpm0k2gSZXF/fxnj78v6+/EP4ULPb6H0O21Qad18yUSj5jJelRgrPxNDPFM8
Nc6FJeu8eYAjha0kxVjrfzuVld/DoIOcblfzkcwX6mZMKNulzZP9fIahYJVIJup5OY2lF+UutCID
gM9YkT4at+YrtABTvoynaAVPbwmAb/5MG5K4NX9kB/gQrTWPIcgjOZdPq726w8ubQSb4m+m582Kx
FIaW+uDQLC5/3hoK5Qc2V5uNTkMZP+fze9+fh1VIQ77AoQtQe9RwCUAhUFMoLj8BpdmrP7941aCp
QMx20Mu8cLWKsgV3s83J4azrrK0H5vVHxJtN7SIYkqx1TBS2HUNvOC7AfTfd1s2cslYmVOu/JIQ6
mOCFW8vGDUh4DhqouUp7IZ60EM4MarLjPLcmLG4oYP+xfOi6p7K4Z3pzPyqc73dr9YdX/N59R8vJ
8s6I78ofgGyVXuRykZQuITo4YsCsJQNn3F4JZz+/VBPQr890eZD8K4MnakKhUur+L/9SazqAcv6b
DACPH9HNLTwykZ4+qBiXmT5Gx8K/HIT8IxsMy3i/MvTf9xJGcBDaQa8/fiuDIpXblcEJAjagT77n
Treb7v1nMyV/rL+h9ch/clxX4b7ZlBa/0DZVvitPHBE9fhbElOKaPkVfKfTKfLVDSdjo/+CNMxYS
ZVze/uMBoq9bjdp48tTFeQBhN7CpY4E7SSuVKGh4dFiJ+u5JvJisOdILhCt4vD5okLOJjubYQnxv
+PulLqALUyugMDrYM1VzvEQ0KvUmuBfmCVwfVX/+BGaCPC775kAaNd1SnFiABOxMUhPNkY1kIgBH
oTEhrJAgA9kbK9uThEXV6OBUe5Ymmg6x1A3jg8Ez9uks/P3s7rNsGn0tRLsBs8ySaLgNpT0tc0cI
5mILDOo+ntI1n0FW44TiU1Eu7n2m7VhbyS15nB+YRgohxEg0UjT3rIWkHJNUcpEBhI2wNRUolS7o
vKEmnRcJ0PZauN71RaOwWDi87OnCh+bRcug6sGFkG+QiPhTrN7BBnnkAQPZzvYTTTj/v/fI7tOXi
RuDse5P4h+4MOt3vBVgafBjC8jwXzWNDcHStl0enYIMXb1EcLAiCj8g0W05z3esuYbA8zCCKNhap
GRMptAVX+jcfH2skdcCsWq47a+udSS+xwHgAXLFuJn7l6j9jM9Zc8eGUl7SFmVMFBVoUnj03OMo3
h5er/EVHYLnxryvzs8l7CS+Xt2+7V7S1Feizl5+E3UoEXaC4Yodc49UgdAXypJQE95ju7GSa36/I
9hdAQUXHB5+YLGvUHz0OnpRP7UqVnGL9koamTfV2gzoo8PWV0xFI+kpOFIt7KpLpwBi5I5LUuZl+
zAstAqg5nsw4wqTwUum00oiumxjTGExZdNTtBf0MAkEr4GW7ngClUShybmjnK6f9bNc9NaiJ5F8A
8Y1Ge9DwufkF9BX8aN79jlGKM5hOtcJ06Pc/l86TjeuEzM21prhEhUB/H+ynDmOxQPv001zuDJg1
7DVBQekaCY7TCiudjlLyAJXFruoj94aUUOGIx8GuiJc1BiPBU8+G3I8bWYB8VuNsA5sC0tDkpiqQ
J2unOOzZs+UZiWFURBmiyXvL5Rika0qA16jvtqql4eRwRUczKQHWH3sUBPzMC4YlSSpFAI4e+rd+
sto0o9KO9K94O13KaVOuP7pyuSS3pnZIkhs9gGr/emVWLpGsTBG9v4CPm4YxBh+QbgGLw2x+DlA8
VgCYqWSesdieXqXBravIE+kOB8/Qtsm/RY+yVbYdLmqMnZUleINpow3YRaF5g4r9XTJ0vFN/Npuh
ZdofzJ9VWG2Z7zHUd4XWbzVJbBmJTVpNQ7NsoqSPpOVhcJt0mTNTL7wlP5vBVJmWKTn/dU/v8hai
Smr7/eDhFYdYRTSk5owiZCcijFxcelpOc8PhR/4Yy+TVJ+LYg9RjZ7dKnlw7xnBEYYU7EX2a6i2x
cG1UvWSSSk8HQFgFgcrhT5w5Mv4CAlSFYRFJgBKQ/VdxHyBwOaVtsWKbGVBl+PtGZZYRQvsiBCD0
M6D11RdgZD3mH73L7KT/y+ceXzIreDqVrd3nw61mWaf1o/bHJCODu3fka3V+k1x/mcPcz4tJbm+U
4JgD/FYE2avWbAi4R7qp3HHTeyWH84CVWvjw4K9+jIrTMEIbQqqKUdXz/m9PmZPHVT90eT79y2fp
teOMzgy0D22ZSpEAFW/Dmn55JGrK5vtW6HBcHv2q2y2M+r39up0OdxdgTv+L7KF75GMDGUeZKfsj
qdYQRnmdhmCnS3ulEf51potQdE7ZuopfAQXDzC2zCKK+TOxmoSH/NcOUJCJhp4BIrN/1suWFCDJM
rfFRmOxmGMT1oZuCcec/uLLkN/+ujDdpTVhrPlkbgheDQ2JttOZ0s6STlk89g5QAuzfqRl+jb5Ip
dzlQ4hGt+anLT0NukvOra4KAVtw78fWafsVxPnm2KkviviXXw16B3+1NZ4KVnC+eoVWOVVTef8Ve
iqCWPk1LQ7EGVe7Ph6QqIBFvO746mDXI9aWK7vD97L2sIbnMFlzGUrc2jFzda4GMcBL4Fc2vC8Y4
1Ax1b7JZcIkRp/q5seWVw6lair+GFDWXa/ml4JouMu+aFLNObVlEFvRciGazwCTXELtwWaZvR85B
tlBcZ4gtwVIuStSVX+4cW95TNG20xxfB8iSYcDAW5pzUhtSN26TG3IDzKE1k3xFIoFmrorxhZliP
8jn7inTQ7bvR+HvTJHLFMESF4lHc/DZ8hJbSlOYASwU66qNvGg/n0BTe5nK1CU6dnkajQkR8c6YA
UEAFYKm7gJnOb2P5ilT2kjhkDjunPoSSMwgWKVmhr2CSRYLznwLyBLxnEUvdM3QDb0dl7j8tfUeU
v2ztqLu+6FIQ+ONbeuAh+eXu7KzIvUyfuQhqC+InbJzBSivWO9JAoZuXLTb/xDrDWmybcPkanopM
iVzmNicD17K+DPicT2cBhKemego4asBmHvznALgXfhXzjTJS4M96DtIdFadh/zhTTirEql4jMU4e
hCUR0ZF13eyafvLYnzChrkHkO2xqOg20QHpJnxuHDvvhMJAd+LNWQGlX3zCrMwl/wPiknu1Lzd1H
FAeNghwE7SiMvJqewguF/Dmz/lBVIpF3Af2vtO+tuxflF8NHi+AnHEqAIG8haHd5WkPUTmRYRGtP
9up/smsfO7opvgDjj+IUGfwLr/wBLGdY5AETeJtqUKxSRgS1Weprh0deLan2fcRX8k7SCh3ab+ji
f0dHp8dqiPZeTvCt85O02FW1hrCG+F1zcQuP7W/iukptSMfsf4tB4sn/tL2HTFFsDFuXhI/azUZn
yGG4Cg7g/yUhjtQ5EJd0fzcBf84ZEYepJMNByY+BFm+W+Lcw3nxLZ05CgOYKuWSEu9CYTY9ALKJA
NeY9ZW/UXTjZpKL5kk84qCgTPSeLtrLehN+/nXoXlih2vnMHPPWb8M+ZVKJIrHq/15fsmtz3UNIn
RECE6oVXY46ts4LwNrl2Mv3EvPwesCcCp22cq2np9YE9KCkBy9FCG4HApuvEmSarsIe1GtjOpjs8
D4JzD5kAKFB1vkFvlxSDqz+Ab+pXtlIv6f/3xIYZZRf8f7gFzvNcITWHl47h6tdzegi7QK+49gVF
P8wH05JFwDCcMwymc8CKw/g0RZZ+HsdB27ehJW4+PZlt9jYq+9143ou+SmgZA3aq38A0k5I/wDKU
xLYHlq3iSpePhswEtbqiTgBoLUNTIe5tkeRA53ptVPZvf3Y3Fvjzqjuqatvr+2BI8TgssAxPfKTM
J24iPwpuvIu1LZIPSMzBiuA2NEY44zopbYxcPTL259I7igCDmD+bWRzH3sSIK2VmFHqQS7fR3RH9
jeed4G/J7Yt/iMr2FX8OSQULLKvcb0IoFGWYP9V+qwInKFrJF/vRkrhqXj/9w9TRNGvPG6seYb4K
OBWEuuuc3xUtswFRoupVe0yMuZcjJW+Dm+/CSkVlym2Wv6rBM/wvJCubLq+3dveccygHkrGOJ0XB
fMWBM9j07fd16qhpEeh9FYc9oh4kzgBZDy4xabPVF1CHujjkGAaAjlhcQ5KtJBIIV09u+jTuXCAq
kcZehkPVgd1BMMfRX/UIZgpTig8SxcbIjdp96Yy/fiDAT/GGM+R9rXfYDq1uQEfGPHkl+HcE3ZfW
aJ/toU8vVpVsl0uMun5/uYLuhYr6VqXV+jzf/W1Eqi+ifM2rCEWH2GzKxDQjwiHiHQa5wm4N+iGf
08W4OIy3bhnFt78YjKSeu9meUEwdZYkPoj4MDPhTuU5NTrxIFNO3Ri6SwhSo4TKEBbjGCvnqrJGh
JnCYp7+uQMnFb8ZK+lGXAPNCWHKNg3uzNy1aj3KRJ1nlHbVUYI00gyOR8ZngT9NWw12c2SN2OEBJ
YJUPO52Ixmejk9kaLpHvjBVL2fCEkX4xD3KBP45PvxLyr446uiDSGkTC4pgrgpd90btOLFjP8f89
JFzzOMeSOSyMW9Fi7nZ17HbXWtndGNUCAqwsU6r/0B/NIr7+OvwJUQXHwBb6GmjXhqm/N5AABxZM
XlaMug9JxZACW+FmsDsJ5UHB8YuaF+JjyPFnYQI3z82in58pp3J2WcwNdyJ9d5tQS41AWoQBJg5w
7Bl/VsfhbUA5zDYFnCinXh5/jnEPcYnVHRzUl85KTA30xA7377dhW0ANFOP8hTbAHuOItY0nEW+G
ft1LxKXk/4sgabihsbx8Ggcjuk5b75zUhBuz9FVqSyN27vp8CCf73I7Zq8tl+2B2xOTOC85z+rJt
G0IRBgz3EpGO87SKUzsiUVAUk5hKP5vvHgq/GpcXRVWfLpWOXBgFqdr0GbcySPhdxLLw9Xd/t6Ps
EuxWGmVTyjtbzIMRxKhqBGnIBE7YNVXLoWuyarKN+TM1n/b5Uvh1hGM1BUBHzqinVyvKGtx/47v4
R3EAGMHLIPrs9W1UHurHBTALILCB3ItLVKel4Fo0WWXyKFGkcRTCpqCRa4FjUBNaWDJT/OYHqW1M
QBPGhd7FrbKetDSfbiWGPSMS0DQUCg3uqMjLxjl/lz3UzrsON1ZwsPRLH1sYUoBc9tog7v2Lwq21
WLJQ6T5i+bZgvETGuaZ1VyiYOcedN9BRUUtxiMgsqk59a/IwdzNBl9rUTxgrHSAPGlcWtR8o6xgC
+m71ElLu+YwLe8q4/LJqEqgNMlEBpchT5DuK2maGB5SSwReSlzoX68pXYqQWPG9AyS94es4sUUIu
n5T6emf3UvsLFpcCZM4iAmjTBDzdFG5swSu716p/sSucuLNCBEgFQEcExjMcZ/MwD+OvmuBDdNdb
89DyZhybUYHxJE8/FpGQmUuyIQIOIcAS7ZNVB2N+40UkANwsqMrcwV/JopgQ+g4R9mFpSfv4TaIn
CMaND8ghFICn5Ms4U59+VxiI5oK2T8WGnMKTJYqbBZ6HSMmx6GqW3+RwGnaNnvxRdHnBm5YSIAGg
05O4M8zo7QtrD8b96vlkrMY+/ySZRET8RIndwqnUSrVRvuGdwj4HIM7ncOPJIMbhAcNMTAUm0KS9
gLT/IJnvfuTrHlg///cRzsplPUfxNKZafZ4nhorDyNygN2yjnolz6EB6X3panG1z7Roun+AJ9BtD
QL8cYlGE2usuxWfjMqAT3/3X/f2ZRw0679zOgyn3oxxCJHQgBKzGhraktrdW3Dt5DpBQ/rcAR+Cm
sfWWAbwBRBSuNYen6GOCYjGaOVNzkgsUvwQ1hVrblrc4PBbG9loyQN3p1ndfQUgzpjVKBCW/hmoo
wfyeIArRcHhPPLRZ7OPMGtrv/4bJxq84mb7R0LbCh7e/G0Ugp5YZu3od4LgOcuKHy1XXiKJy5bfa
SLwVIekav0ujrACyMIvTV6VCw2V87q/JWFrJXHsi0hV2M1rLL0V26IIM84xVD3MadhC/vJkF1krS
nrG4E8PREGdrBNgDIORDQOYbfrO74m6Tgb1VQ1oip65lWUigj4gPNY6QXqecOBr3inVcjkikC61d
Qfq78wYND92KJ+afJJ2FjP63STSInP5okoDsnOV1AgdFLZufWI6qgjLZYKUG6uGPhcE9zlcx8bXj
xDhD8Cm+6rLVvPq3GQvXGoGYzsArS6PSw084j9dIjAB17xtwOtXZQi0+vE1EEnKQ08Ao4Sj9Opae
E4OW43uKfQXrbodp0S/tbT/ivg3qfYbKWAQbzJQRNaIOy0D76CF3goKJ+D1eVCrLBY48e8G5F6/9
tbtaXCWFVMz0/Hu7Mpt386isumpuHqhpjyG3p7TwuGUp5njOCW2ak29eeyZQ9Pw7aQnJlvrUHIrb
/0yLTSRPmR8zr5GhOmdKGyI2KULICciJZx0wMyfVwTGXf1nA3Pj/Ww9uoKhQq6jjR3xzyu1gn2Db
A1pNdQmM4CRhZMnHU/MqSr1aQK+gyHxso31fNRda6skLZ4Z4ITwIrSHxj/zJ4os8lC8Fib02UnJG
gbF9reoY13FaHeCqqXgz4Dc4L2+e/MsEABEyLpNDnlCG+4IxNkTwfPUkhlRNX3l4Bp2y5ikX9U92
vUyuAybJQ4mghYdh1UIbFYbcPUJLw5Fe/3ooTfBTK02CfY+QRgJ2KozqwciWliVpoNFOc1SYqIhW
SbsEOnYNu1t3TeIY3BHOv+I7XuIBGssJ6sxfczMuLwUUNVDGTwFI5Y/XaUoHfkLwNd+UulfRUmcr
U8qJXVbGum78LdWOAkYh5no8UgPaucLZyHjOLRLkC+VbdcLfwSs63KTjIDgrV4a3uRijWW2D3L7v
pkEmCXxcFVM11eEprUpGKwVC12a3CYL8b2/IqulZy1oTd1OUgbBfM/BXTWhOIwZ5rrQaGvNYdgki
+8WchZpQ4pLkM0ixYXvvfPtYHpYDUhJtkpy8x9P2fERxdDJeqfO9vRW85Tgep91BeENOjvNEewJ1
R9vNcExWWHA+noVG6O2+ybA2wMmqMlvjVW/cnhuP4fzFy5TgtAX3LfumPNDx9BsFoSb5G2ke8q49
96kKaMVAV0Z+sk0nWIG6XdlMUAihFL9UB2SN23b+LaloQSvQwpkoADlYwEK9XIF7tHiLgu4rINEd
uW3gzZmGxc0wjFlsHyt7pKUIv3xA7xch9LVHAeQ5ajqDTxW2GyCE9rfzTAxH5331SbUz8dt6em/U
Nnvc5+g8juxLtFDkK0HxR5KUOEjSOFVLVPI/LJ1geTMBaDHZmIpVlhcIpyiLEA4utHBPbVJq9WRV
l4RHz160HFs2G27fI+P8J/RuakhU0Pf9TOvmXN8lrcZsx//O8Dj+QyHhjIDsRy9aIQ5NsQ3jfOQw
hJAfmVeyEnsgk4hEHUuPZ8by9y+QR+S8mmJb+TNFTB35O8dw9UT/tYfTIOuf8K3xwd5bQzU0Qyk2
Wx9JcTiu9YWZP5wv4OsRpHIgWl7/jUGKvNV/w8A2Yg81tFosFGBPan+r7paPzmesKG91kPTpzjje
nNdK2Xib/hkJulSK+wbP9M8klhmTOVE0w81ZFUWtQ4SbjdH9eSHCEe7kaiq8s7w142mLgS63zkiU
Q32U0Pst01A/OelwovjhvTPpeNa6+tNES2mNHUE7cuN6yTIGHjh8aFmxRDMiefM2g9F098jWiekk
aeLZ3BEVoer835EJ4SDo9yWXNxdkQdQFZGkaPY233GJSLTotYEsCOBoe08wa9jFI9ppagcqzgaLJ
8vkaAjg2aauEsDdyMAv+oGBl9xtaRzO29BTnPfznyhZ9feABp9uefSdx3pFwmmwjK+YlrkcBqFUs
nhbiYHlDwMINzpkVdi6XTJmQP9PK8Msq1arQuvTof3XHKTyR2gpin61xtet0l5cgGaAeNk5H3bwn
Kcy6l99Zep0UG5TfJqACdH9AAFcBh3NAHHzcG2QXmzMs4/jC/C4Jc6LtNs30lfRQZVNpF9BshMVC
HaaXQ6BOjqrEVvywOhls6BuvX9kWOvadvXz+TjKKF9g2eOOXnpCHXZ08kcm61uAtBeJf2s+y6Tzt
ImYWH9QWaEj2UXB6Cv8CZEUhlPBhhPp6e9WR3TfjoKketfA7MlypwB0kNJvIFQF3kxBR7j56iBpG
1sBq8qwbQlY/5S41+Fwv7IJEO/SULejNmiZBvN4fZ5ihvmvEp+Ivmwbj1yHm3GscVrOSpnjS9B2e
feyXvXS6ouKyZgwE4Fh56j6zTUPabklqvMCVrmRxKWmgGOWo6WfzO0PXZDNn/wZiT38T16dCx+Y8
qLHEBbumIje2CeW0AUbKK1KVZmx0G6O/68Say6STMLbVlCkMmhw+JJsC06D2C4JDYg7TfSCWc3kS
if5rCz4Ie2SwLRszOdzRMGn+xhMsmr3FxJw9QzIzQYdCVu7oNQ2XsVsO9aR5/TaezUjZaY/3ecAo
tZknM87XrIunJkoS5J1fmGvNbS++LhCqPkwNbG58tLbplSTuqzgKwI+vCJG1Mt7iU2fmLKgM5KQk
8g1EfpaWG9uOVjdYjJxonMfV2kKuG7WYHrjoDPGzCCNeyvpOXDdzHCeUGjR1TYEcxV5FibFZnBQH
5Xs2vL8xL+BAcas2mFBEeiPcZ2ucvnf0hASblCHfQcQ2+33kyap4uCDsCIbmpRdH1+lCan6ECARo
PU5qCss9iYuXnWgmPh2bHWlWydoIDmTPvtjB579VIqG3g1WB+kawaPIvQZ+sHbmsyyXLLf+Sgi5T
2D5ZakVY8OXITE3re6qTJKuKhSkuiWuVSG9SfMv2jad6PECaq1YUb/8DHT1JQefcEBSm7yQ6n4kF
XQPrCCph/WKJdPJgPsYKOJ1BS7SLSdQlc/Trvlc7UTmqucAcu00WKxB+o0hUuIIME2Bv+WTV2LzD
uuNQjUQnL9r6+LlF46EolQ4DuO05BZHXP+HEs88+zaYxRtTR5xkBMh9C5cy8wx+Y9bvSEfS+GIB7
qWg3pV62zljF0qFtmkZ/ewvCb3ViSucJvYZthyvHSJ6rDZRfOLousIo0TejcUBVru+ma7Ss7uSLe
wrZIqWMJrF9+GnFGfwV+1iiEVFoybMBK6l6yn4CVRqHoK+2IR6xZLLXZ1IsedaeETWiY4xyf1uHe
HSWM6KxC5eUWE1S4QdH6ENaZSD6f7jcUaJY49k4O3iobWr0IGC+xF1LybEnK1Xo5jRfNGKexseex
pM9aOIY9ZL0wMgdctpuJTHk5sPHU3a43EUw30jz/vbBK7IIgM11erN7eog79WCUt0Rvt05tyXmna
svSQR4PcFqCYl0MbqqVjcE0wfUE9NqvgyF5q7/Q0fv4pv9oV0W2uU5hBf4CEHNUFUvvojNXB2V7o
au+PTYeTxBi6jB+4DBw7MsoDWX6/rQo/uxWUUg7kSF5B9lEQKHA6E9Hs/POrL06ZoutDg894ZfHJ
CLTqYj6MOs6h6SOcBRyt0c4q9cl49lcCARc9isUSzkPAEKvHiL01OGYhh/FXj+C+P1ngf3l29HOp
7ZvkmZ7tq3hl7ePzNct6Gw19JQ7OqQPHzsPcJjjG5CMCVFFm4l6T/CMUbPnkmC3i8qoMDO0C6F1d
+YZcIfV5QTXbuJn7Gr7qj8C5VrAplyDIyqDT401WVeZRnKWx5undqqGpKhSrIo8EWNv/KS4TuclE
g143bd+uuqcz3PF95sXDcRCc2NZkjbEA0GdUUgyxl7OHX0LYRbeWQjWC5wnGbh6VpxB+ORN/OqN/
A50XOM5MNAOgC6fNYZrNdnCnTsbFQEbwCEVfuQAkOMIR51CNiyRJgJqbGag2Wo1NJp37TAho1W0/
VyaHa9quFPLkBFJ7vT0+dDxDwbfKw4L+RIwPbfIYjhd4CD0SWwzVgVWDgZ8BY9gfeX9L7fElZgm7
sPmMhzml08Wc8hEMdOv0rcR66xZNYYRbmC/bnculdy1A9MbRDG5hTrMgg4Y0qfmg5lpvj8JRE8Zy
eN2RHf3Gr4BSqZSU/8R++rKUHDCJWWAAWkacUpK/5L6EGA1PyYPwvCbAprtHleTMLQ9woOJ0LU88
LQScYZbaqcgeqgHzQ5XJooTLq1oeGW6X1OmX0JFtNmdSBH6uR7RCO9f/vnpyUUl2HXjZuWo9vge5
zladlHuGAd9cOruiNScTAq+nNTaPtKhKsWzPOp8LY2v4p/CJhs43J6ufGp92JtK0vZ/zEJ35bK+9
ZgF/h3dPU0x/0sPWVlqB7Aqr9KAxyVei2LkCOXn/MNCZNvGchbkaY8Yyt8Ny5HOPuSYzThBQEUtd
cK4qxhMf3MRozSc1+cWU9QjeMc22w5P2zfEm5Oz2dIHzf+pyNXtj3FtJI6IOi8cd1/v1lKoeYbzw
WWEiDNbaLkKImyUDyxSUrCKUciCI4pMLgtJgAh0JPi0JhWmYY6OOAU9ojXnBg0fsjjWkwcIodhq8
aFsJKeVBS+76Pgi/jg/VNtNcnLiu/1zAtQgkG1XDA6tFEBCee3J7PYuNKneW1exYvolL1GItpUuN
dpQZswaVSq07esUiJq/CtSWUY1hFR3gtHtBDtGR37t6VvjCgn/d9uQKDDpPgx6oRZDhZbzktYykK
oPnMNKMtw4Ih8Ti4sdCelnMv17xKDrSXslv9hcdALbBRM7Pbj6iRKm2MQ1qpTDFomfyjH7HLnRo3
/0wXJYOj39PDUpwddG55zr+QZasSt/muOfI2cwGLJFMQY1MI3U7BoWYqkPNCm0G7PTXyjm95rht2
7x+5yMMMxNRRlFpAooKF+K9rXJ4hTVWe35ShQDsYJPMotLJyvPZlG0PpgQstVibLwfx6vfKV8Ald
D3jvgndkgK1P43hQP36LKhdcBZFWd32+Rl8FblWElz0aJzIji7rRYkxLM6XwPUQLwpsQvry/thPO
7rP/OEpYST+WAUqWsB8A+7zXbUoQiM8NjGUupuFoobnnr+KVEKqG9RGHk7436iehkuPuJIdrURSW
gXIANMldvW+y0TDNTOmUeHVHrXd8wUB8pwgYaaAt4FKsqhXw6V6alaYNJEh7ncW8vNBnhrU5UA+K
+OhkSaErc3BBvNGSbHdz6kaJdDUvpq9FufabLeAknva9f4GJKajpJ3AHbp1IbuzftI1HvXeVSnap
mUiRRqFAQvGHYAynu0IEg4Q0jo6rM6ngF4D8IusllX6Y/H00dHXGAPLHL/v7W8uJj6M21sP1Ed5v
oGp89peapcAKJNd6DQKmNuc5lqLjTDIBWjLJI/ZI614szT/qZ5iKMhMJktg81kjGvzO3fJzXz4hH
A3pNfp+G+S03KGh4K1V1SzDyOifDRgBXOZkMAHxXRaRMp1z+tKUfDBZGdoXNqepGJwGedLUlODsI
aLDZycDVc3a4EkCJUd2GPQOCKxcV38BcPAWDc0YB3lfM1HTTE6PRmzZIDfCbN581hVfzxI+F4Suv
M8fAL71M/lNG8uWLhdRkHxpzaljzh4KWeIPm0ztPpxkFUPNn8cM2trqdglsJ4ZDLAhK7XLXpNWKF
rDWhCZX/kwFGM96xsw8/jQ+vMhbFhOObIWsXUGdGzjuleXzixFG2z2v3YowQBbbf26LbsbsIDg0r
hedECme1ggUX7/RdMhVeHlYYBd9iOzQaxqs/II2ZI7rrresdLj1rUGB6L+f47Yt8s+wh0uPWbVRM
hHJlS9+hB3L6uko3FzB+7nk1uqDj9grMe7o1dKVlIX0gamsDj7eIk+x3cGsYnbiXRzmkPkYqOlRP
S67aftEjM7+Eo6Ac1m0vdgcmDXW5U5bal66tZHgV8RDd9GJaRWaR7F81ls9ZNj3fna2LaEryAU6/
L0bLXqtiEcGlNnlj9pgFiCByxrhhhcwbMzA4gva1hHsZtyCMJDj/ZCPVXgN3IIFLqv8FXWf7lNDu
XZCvJUKHApbGvvKH2bqk8aVe3gHYq8sBBhczKR/tpP/Cwi9xWoUrOM3M+qWmHG9/h8rfLwkyQEbu
1ZiKzs0P/X6oYp3u9KlTfaVK1hElgaEkwKbfk4de4h5k26/mS1Ak8T+ymUP9hE/JvInwVNL2WP6/
2nBkRfWUYeOAvsyCE87MtLoHTmzNjlGIx0xvtv2vbF9tS3gI8zNwqcfy2Wr+AND2CXLO76gl8ib5
OmGiGnMBp/3POT94yjSycKt6l4yN0QNLR07GFLlEpPqgdIVRP9VUSyk9f+r3FX7mvcGQvgHvtBmK
stuecvXCyp5eZ7r5TLpgB2p+67UW3pwTeE7EMsLfvozbjrCuQvhgipo81Mo7A30nfZKVzoDH4cbj
/ck+XRtTYuWLUrJTLR4laFOkkwXeZAFOrrMY6sbO0FclnWJalgE9kCH6MBiOm54MXcSY0w7Nr7x6
XJlnHL7jDBEmo57CDiofEPH5PEXa2A1E/G7NzvXgkpSqRO+iXqJw5QBPKGhutVRDjvD2Ob7NZ3F0
aCclRJAQp6HnAqBffXf8RySl/kN0+V6BparFhyzm7hZRkntr05ATAPqpXJJCGSNGU+FSBta/vrCP
XugMLs8CGV5h4Hvu8EebP6sfnJztK05jREUqFDU2z+krrs30geCNSa+Xxl48DgBpE3PhRyM4enF8
vh0jfn4C3hytLOJhZQVF3kcKld1XC4Wbba8y0NsZXcrCxvSoqiQLwNzroxfnjuB26B0d9/kFj09w
dsr/mS95cy4CTGhrLepLvwWBreOksUiaQ40Q8W4s6cBvZ3XB/FAe1Kf5+oTfsXGqgXTJV37uO6Bd
BfUtXIxsuf20UuJ9jyGeO8ZulWfUS/prrMAhWtkBdmqENmWy71pY0IqgDKG+GR0XaTyYKoenCJss
4nmcG8QGLta430nuLMMKz/DazMzNtKDC8ttqU8YL87KiQvQvbQJ0l3TXY6Y2aQt5KAXVyi4g5spK
L8te8O19lqiAijS7hqa8e5V2WpyUFGIXRUAxzvMnNBFUgqZR8Ehn1yF+/qInlnghhRuQRjDNE7M/
Ws0y+INLYON8VGRvu1pv/gYiv/CODKffi3hoTu9dykP4Ve+mP0tbnVcEZhd3Urp2TSh4rXSVmtEq
TyLc1Wn0vEHm1U5gVI3tN9pYx0vvFHfUg1ISGTZdZtcoc5bt1HnMhj3AuQoizq+1A4kIVDu4wZf8
9jvFNBsJ7FbWv8NrY56x2xz+McSIEN+5PnKDYiks77UTT09kIkrcL8pzGc8nCAUxw00ygHGmoSN3
vKbqSHFZbXccTbri08VXarDHegxpIDwPdryIFfLzVh12bGPocYIFIKU7jfB9SG4rzoyjT7RlfZIm
vIXlnIzknl1RzPCpUvjTgpP3VICBRAy9EiedX6/A6Qgr6kSHbrtIlZbwkoz6dxSO89GN8vDrZ/on
cBeACyy5H9hPSqAICMJqK6wpG6x1Rr5DCm3bTA5ZNFFKz4FYx6jnSw48mnS4bhd2Mw51ir4ym155
RppMFKsMs5hT9WsnthisJfmgTVbDBD1Yg4o2u0pN1W8B0iK+A8z6CCLfVLuqBOV3t/qIWLov5ACf
57sqLj5FDOfQSGXF/3ZVY4Bz9XPDDPkE4JEYfemHDvz5ZgarJJLhOh0JNeuoPiUQdIHJMb3To2WK
JTIAvhTYyqTYcujywfmLeqdohzLka1m93mJO4Z3JaYMCfzmSnxz7IX2VZxftma5t/HLGt595fr2w
I4r62xUQtdV8bk629Bp27ETZ7NGNIX1Ti1LPYULQugdjsCraaI5uJtqF8CRwnVPWple3OFJ3DuJv
RFJSpJEVw+NQPk4K0CxXI17M55BuuLgKh6B9qM787/jL14KrafjtiO/9ruRO1+hbElSW4P3zGrV0
GSgA8A+WyS2lUuQ3SBNBzp9fBUTTD2kp/jQTYfCgefCkYHq37u5b6AYzwMRVYVmM7BfHP2RKzmuQ
Yn5MLB1uksRyRx8cY/2Z/YvK/Zgiv850Ca48aIFwxT7IDtvlCTOW4sCOH7dXAO5TivfNzgjj8o0z
dOc5OSnLcwN9ELimIUd/dLMr6dalMaBxSiUBmFOAlOobwkOQm+jIkvpaBWF+NN7b1TGVS+BLF7Zj
4SutXZq/PjIO0UDTh0VlpGCLSIaubrpH+y2fDd0l+Zz/JwrcmYbLBMTo3f5xLHmxW6xxCc8V4vQq
Tuzb23tAcIPAwuWsHFXxzi+tMO/UViGkxP4q09pFfF4/LygM/ickVRzH/QMRmSXd8iGMNhtgcnMK
+C5CZiQOqMEm5Z1RBnL4i8KIydNcecti2UQ9EIPk53eF+YP0rUYlRw209jVaCJSzWixMvyaMQabz
6UaatEIloVuLY+ejLJPiHJPXVjMILPmCTuCS6UAuIhSlf5f7+FDPahakVtLL2JWYy9oLFNa3juca
vNmPUsaU6rgea5fJzyA/uQPV1vOAA8bzLSgHPBuGBULjMVIDgeVpqvX/fpqUh/0x6uRWMWRYWQwJ
Fm6WVVxLK0RgmZpNlBEqG+ugsRbm/ocIBkjAPKDFxKpxBxWosMuz9u6WCU+VBLfUO3opAkWFmHZ1
UPO/2JS/TwCZ/NIwxnKJg/Jwvk/nH8vwcu/ma54yPxQrHiXOJvODcDo+uiyFbKIACbroCPhBOC7d
0JvYB44FcqFgJjVcBu6O0lKB3J4hKWQQpF7J3gTXLFbW+mWt/kyjCVQXW3uNNH/ho2lqduIJocKS
gG9p/s9WrkhrJjJI5nYIh5U2II3xI0131ka8adKiyvCbAGs1TiAbq/Hn50aLxwYBnh24eyautHYI
nkaAAwUVpDGxFLP+YK1ui7n6ichW02/KM2ceyFxt7EQbbrqiyIBJwVkJ8gc/142ZhlKUy0IwtCCn
ZuGtow2OXxx/IUa/MpgbufeDRJwmO3MWmy5WIyNd2vNF0SbMF7fzdfhFTNd+j4ZMrXTq0ovH5iBP
W34oGSoTjgfd7aDnEK47aiYJz3TFZHXG/loiJv/QnxMpv7Su9IqM/fd1p1bPJLx2VOv2UEck0UeO
OvadIgfeT6mFpxmZ+NV9o1wBHSo91YIuWvHmQbW/imcziQMLY2xXSrrIMBtsBWSvzOv22K9bHjEM
IO2wz4tVplgcx3tvtLdwybSEDGxzwPROhZ9Bk1gdWiLnYeajxfBESbFoRFbcNyaKDQQEqG3rkrNl
iYCpi20kRMX0Nwj5AlLOh0Qx7/Etd8zuJyQjdOwLJFGKSc7ZPsGVUwF5tyWQ9ltG+LyM2DEvUnN1
dCI2S5ADAddfbPBG4sRXgFefCoQxs8ZoO/mwEx6O0ipGCJH1Kryivsxeb7btyLK5n4BLXUfnR4Bg
DZ9zP0yICdmvs1D/iSi1N+DNXCli7s86KjGGABlkKKgl+30oczmiJF+Yp4jtNezVFaQ5JD/IgZH3
FbZ88aAGEfxBF55X9YMXLSxuFgxiMPAvoC4Z9K++NPaytUx4+77IqoVlQk9uVYb5HmGG3ou9lxl+
qb3m7FfhoSGaWph2YTWgpQVo6EZQcD1VDLm9b/K5zBKX/8kCsZ+abx0DeWQGXtRjsf5TLneQLOkf
H2cyaObd4saJzBySOig1Bw1zg8laW4dbUG8y8KonYFKeD126jBI7A/CIyOVLMtpKY8hAlEajTxFX
PoiEy33iBVUVDwMYE04ZJOQ3/O7O32QFIHEPYPYtjJalMd2CrsGI1j7ppHYVk9zVR7Rhx3UnYMPT
k5x6lOMm7qs2daQco+FvYFseD4+UC1DenCxx3UlDpJeAFvZ5PNvsbvah2GUdGdaqPGO/2/NKWizR
hkNJNSWub+a55VESx6d3PAXkmgtX8GVP6K+g/HOtIqtcgv/SR3Q7FJwCeGN7wUh0RDLeDFaziudi
juwAKZdGyYA0gCfuxD/hkU4q9HQ1bKLixseZy5D9LZ4OsZDvKCYnP/q7fXLEn/M3hJACksbtMDYp
UzfW7DHpwt+p+7ZSj8cYwmYMAMSP1jiAa7hdVdaBQS30O+0GELwJidFt9gtolZ5Dnuf594QjxVDT
SriAFUIzxRBnNTbWZuMMV7gFVPyjFsVLXcK0R7hZiGf6UPlmsW+QWYu3iAzMc0p5k2A0iOaR8Vd9
oEN9godXrA3+HYnu8uWpHFM1tu9lQX7e61e6H3rqJKO22Pqy6Mw19TAMO2Cp03H6kLSPmC4p7mCD
wp0VOI8xgvMSLH8/TsUHyS95WF5iy/W2fhY4TuDhLqdK3guT4RKSJjz4t7IFvlBV2Hjkes6ap3BO
5XfwPsxRlScpBZqwn2aPHWIqyG7XDh+BKtEQoiqRwJFNEpzBOEsS4/bROC72ypUtNj7opu/xUTSN
JboQZeuGZT5CahaCkFKGcOtRogFsj0uM/FCpbOuctZ93g6rzJ50TyesNRDr8AJ7fKwpYQTpwQvwF
yw5TR5sV+SryhVd3K1izv6RX/1LjTFcxvKLTqVi0NDFVp6qMVs9nzG1XGaIradVnJDTK4buXoryy
QjE+HbGZmnYtzh2fM8mrDbrQ3imPzakA0C4qVlOjx4vhnGjDVY0u8cn9Lx0jKf782uCzkgvD5l+Y
yyV+/6dGuNRUdPpo4hMAmrcOkseYT/T+7/j/r+ySa8qe+0j/01RrhX4xwBKrUebe+dta7/5xtgxr
20ARWWXIsqjD0ZuVlr/ogk8ylxzyov7pEMMWytEXJnNjA7ARL/Q666qv6xsvoLPaRcgEw09f7AAd
XEjAPHozQYRPGquqrPSKPXDzx1OGc6spo+6EzCwL/A+axQu7tIIdVTQQsKEjNUo7bdR5iRTW1GRV
ND0gx2rOxwO2qkR83nEf1no00UkpfNmGRukEoC78e4eT4ip2srFKlt5fne+PG+Lci2quNwjpiAdx
CFPuanF2VAbz9bdoPrenve4qSKKB1A4lbKnkEay1BeKA+0m3hxztrJKP9nYqyQCz/vwDry/vBXQg
WLSboYJk5UaGf7grLse7Ey5dK7kyNzSL+lkQ0wbqGdD8qS/yr9VXDhGbU/P0njZgTi/bSCAhNobG
+BrVz1U6QWLGeMOlrtRZoSedRWYsqVW3eThnX0USh7fi05KE7WzwqLtg090moYhxq59ciUxcAjzd
9x+4pVhfHrQ0itCixvdpkj8SOfO6PD+4TlR1UCDQigfFNLuH7SqH78DlX9dRGcFE7fDUmnFxEoJV
aFbGdARcMRnl8HZ8oHnBI75GdtMVtX8B5u1pUxULUtdxE8dY9KOF98bMzNkf3BB1lAWh1gGJgXCR
iXIzGWRSdxkABci8YPwqYTJt45atPLSUIwljZ/5t9xZgeyIMd2sdIBDP+Mz7Dw2D9IwbCWr/wput
+jptOxlzAMw/zTV1kXUgkwiGw5krLXMqf4syGD6QL90cB3FTP7fBbFBZb0rElkaXiCIWxq1qx7H8
bkI2l0PWdvvOsQocAYjQRGCWVTv+vNxJlUepjAVoEiyq1rvim9o/He7mxeSmCr/Bc91nX9k3MnLM
PMepNVAriXvQTv2KDzBi7inhQ2fEdFG9FBQzJ/Q8AMxE9ryMxW/+rAUvbyAlFoJVXDO2pPUdPtEw
XEJVj3lX9Zg4YsXdro5v0q+nrLru60J5zyafBEgWq7cEIltxw8FyZgFzAz01gDq4SilaPVDRSNsL
0dV+9fT/p1DiU9jjuB9lzgpSsLg2MvCJUsQIoiYUWPErWpn44vR+fQwFtTeyggOwzseWXo5K8Rey
PfLMWFFp1Ak9SiYnj1I1wLMj/1d/JQOIOs1ecAjxcuarWCw2zHOr0EL2lP3QoPnOqcmEZfzvp3NU
NeEHNC/GgjTeLmjOcaDxt7lMH2lbaTc/UbFcd7C4+QdeYkSQAFz0IXk/w65O1ncqwGysNv1t4ouh
gTvBZ7ZnWbmhyJSYOHG8q3B6ZJSUHps71tRa2jFKgxtEZJEy3VTqSvh7xXPeSe1FMVYmtvHFvX2g
d2PWpgC10kQmbBODwHSPYWsfqUGMMLCKloTacTrfwwk0kZxtdH/Cl3RVPXrEtyItjlSFFUwNAI9L
6ZrQpzMq8cKihBBZjUA27wfgZ75ZOfpDK3giKOhBsqiO7FwDaD6KSzBaCvWoX2+huOVeSxHy6Auq
bIEn8DmDnTPN77wV3mjUFxe1vF9KpGP0TXpO2Hqz3zHDjrgkuJhBsWhyifwRftB6DQaqn9pl2lAP
jThGWyBDXVr45o1AtBV42puEl0+2Ly2tfk5MeitBXXeL+xtlQbXSGSDDPH6LFO6OgFB8dwvgCIcM
dX/GiCHxbq//fy3VOShRwHfP4VWPrmoISv2GehSDZJbrCO3f3oUWurp4xGipU+konbotpsF6KG0Z
KhplAcHpDRrmyOmb5kbUH+GkPZ7qjBFgninu6MmdCTDKW+nOw+hRlfbcKMC4dweJTiXd+gQKtsCs
FJ+H+LsoAmi+c5ExGnRLO1leLPa4zNAw7OWirV+cMBdYh9c0OS2XTHlCWUMY17fHBBHuJJ3biw35
6tiZJKV8ruUXF6HtXgoeGgj00S5WFvY6fqI2Qj7zItxD1vm2e4UMwL910JCwAAHB5/Fj4MIACax7
8+DNJUElvrs3N49yP7/VqQaiIeoMpQGcCmEc8DhBKvxm37biRFBmtUtt2e91KRjgziK9CTtwn3pW
HsaIeZlJ9hcT5x32eYQqKSpWa9yFBVQNLyQKBspRvEDwqyw5wzvxsr+3Ll/0bIsyyr3sT95ZQPMC
maRih53OO2P0nOqAZZUGM2LTJDxcNXoFDBeXsmV8fzDoIhyJRrwrwJJqos+F+4d+pCuevoy8xOvd
NT3tDjbRHBYFOgWXDrQZSmCmaWih1sVvrm/fLs9Rva3MrxB7lh+FVAy3+OLn9ZrBSad3KTghNJcC
KY+7+wvmDTRVT0MAP71ityloVjIfVprRcWSWHlVuifzSePijbdaiH+/jvHDvpIiLilIULPCeLcMK
RoJ3+CVTBv1GdjvqcsInbpAr3qKDvnN4+NB+2hIGzCYQt+V8KJ/IfsOc5eDTHlHFZh8TLMZ5quDa
G8RcJyyR9A1H/lGM6awKPdPqjjBuMGXJoYTns1TKhrp/cUnEJBvqiwrqreZnHY0T9ldzRE7Ax3VI
wafBlzMoKM0Oh5hq5b8OZ1bfvfVlxhJ1X++J4xm2lwESDo9Cl7tQ/ik7WgOuBNJcc2cb/rjMCFtH
C8VuIxK+Mzy0WnVc5XlzlIw5Ur0wuv6Wl3tw0VKSXx5iQK2d7T/cJl7FTQUWotOJfnqe79YHi0yF
JifQDTv3Qeu1i/61d0Hd+aSsYssDtLwsWtLD3E3LljJAVYxmBIS/4o84yeVGGXLF+rxfzn/ZB6A2
PY4FMVSVm3887UsqWIvls6DjVi45lBMnX53OUWsALP0+WRacL6EPIBYt9cRkbwGk9Hyu5SeZSim3
kaK95rCxmDxPKsaFuMRy1ZfACjSdtGroxsp+Hg0/XsV3tayXktCFViWYKpggKMxMFGfD5tHIH0Zr
1OTQYizmaOYCGRyEkMdh7t8VxL3nkvFniPDtsQEwzmGPUp3OSb3qLUoC7xpo4TYc8RuQJhu3Pyai
tJwjQkpAEujV2GN14ai/EqLAYxYNoktTwyJfTRtxEILkwkD+ObsI4upLYtPfDExThX3b+BCo/Qsf
Rs3f5TsOlfB71C6M8feFg4g3hKPOvL3954nJjfQaNxUW7nc5GUMf3ZmFBg8jkZx9kzH+rkj1T++k
IVac/4gUfKUx2dMjI4anVhzUDScXEj/t7OikGlkOTC8AGPg+adxF3VRx/jSfAQfqeX1ClPQO0hwy
+mSrXjb6XXdCZtmv8mYlpb89H6VTda4L7XUO4M0ZILFgmK6NjUzeqO+dDoon1DnvMbGotgXCphF9
Ic7YAk1L0lxcgDKZ+jC5wWNWjy+I4t8jLRBZbHp+6VKXOmLelMFjcbh9Cb1NO8C0W1j4YutySDRh
HWMnuBw/xC8WS/ECy8Bc6p53ukNHJibopNQDhu6MUh11BVpjHyae1y9hwv3eftjHV8gOogm0nEVl
471rvT3VB3BfmgTzJNMq007KGQc3CuHRWA6iVSZNdzlO7i2CMPn7y+0vFCP+XZCIlKxomXYUCloY
LK37Z0vB08LDWuOX63NhHOSt8F9qJoxPQ2QTGNCfJ6oTg29edL9YjIYuYfYp9sUsK/2ZPE02A/ms
243IQTacZ/bhBK3mbZlAf1Ix+A1bYxOo8IT3gC5aUTxrKOWq/lXl0hYNVJBuRkuNDRnLINDRTNEr
VTZwo7V76nmAwTIB2XszyOHZRSeBraCOzBombFJF1pZzGBtI5WuI+iqQCbs3UwQk1wHcP8HuCTvF
Hy06V92rMd3/FFaJphpaVTEx68lFxLlf8JrnLjowwr7SBIf7sVFxQs2FbbMLGjx1y/TnnExg4Mbt
SEEqM8VpU578CB+AjP9PzIkULExY2e//cTCWAfhWOLqJq8B7Yj5pU2VA+CukYbq6AFaFKfAzIitA
ltBQCnMcfeu+GKkW8KvcfxX9Z1fdAF/C8XvXiAiQlpL9XyCQT6UQjuBxHPxMY7259kJBN3gZQWRX
pmUiMToNRNRRkBoOkuIakUZxVAhOsEnCG+iDxfWOcyo6jTLH9hRrIMyRJ//kA9iHuej+4Gk1kVgF
dGIh19ZatvL/VPWtCmmz/OaDT5h4bDYGpPd6rny03L6QV5/W6uGXDf+6vBD0SyGdo+JGJWdjGryO
d1zhP9t3VgDuehIiClRPKlA3YoFZWu+n3zRxGlMvn3TxU/X2/ez/L8trzXTirsyQvFbaOcj7820z
cN9m0dDjsKqLfl4ORQ5AXigm7+wRyVfWHT1ZuuBOI1kxkLVe7yt6AdIpavv/qiydWxRXOcLank6h
1tzbTfO6+rNRG2ZpwbrMQyMqkZUhSqGfHUc0Qnvq5n8ukNJwJnmCW86cEca3yg8/iMbTjMmGkd/5
qlr1k1uUjFiNZw5swQ0AEKzTMvlg+b1MI/PnqDyh0vEQdrYx1qVvfcyuN/7jeGDlpne07tAk7039
jnioeP+ro/Cz5YulswHYxDOk9+CkeP+HKClIpgr1dje/UDmz32Y8nmEMt5lmqotkVuPaVoT9QoZI
txfoh6obiTI2EoMoPHXOEoBR9sRWXgBZWcS4j0XL/5x9rIadDwiZL5sZdzroeUxYRtpthPgRHfw6
Kvb+rUttVSUVZ5mEmvk9QqIH4C764714bopsY8NgHmgpPtS+fuNC43rWklkIBog1KZ4401joOB0+
QhraSHMumhw0yVfjRRag8Af+tMQ+8a/fBDjpk+/vFVl6S2Uu2qZwcxnKIgI4km4m6wGiItHltlxM
pbhVIfnZtMkwuo0rmbpQ5FelL3hX7Iv1my3VfsnJ8trosWIY2dXIKbMnjnDhm1f4lPc/2AGalQ7F
cfXDddnawxjZgFHI1/FJ26Kv6YxTpPQsgEUEbahK9vkkK8A3Y5evvC8o9fttpjznUmr5Ci99hEtb
xlrOGahjDOpkEDK4JCPV/wzNCyNJOLTKcBHPb3NeNAJIXJw0u0bTM9hD7leg2jgXmFP6zN6hoCGL
R8GRNACo83ASmqU8dVy9iY2thH1PAD+bO/AN9IW83o0+fXj3yAo8S/+xA1NnZdCTmfMZ4qrR8YMW
ChUPPui2NDCM1iCFAZzdHibuqg5PAg+99A0hA/IrhNnbCzVzRUMkNizcynW0sZ1xlnGgEvOFTVCD
OsVRTcaPjmAFK/4f4KxWHOsjOStR5whx341tciO5BFY/wYIwG+sAD4Xm5UWDB5rKXRd/e0wMs5ZV
R6z6YVeXxmLxOQ3pHdFsoD7Jtq94KXVjDEih2qJIgGNhqizwMvizJ7gAoQC61+mctwpdI59DHdXK
h3j5J+3IN17lvtL9aF+Xh++KeGnGJhKlauTV6biyZo4kT7FJ/FlFmtMLiZIbKaMMSsK1V9e6mbNf
y0QpL6/V0pajyxn5TDxdXjEbnWm8N5q99QnK9OHWEGRCpuLU5OTvY7nymjDRfIDbiicGN1NXrvav
IydDQ/VA8E4WPK5i7wyxsV5tS8GMmwsTpUHo26z+fhqJGkd0IoSDpr17uDPr/WzV5IQ92RKZLLj3
4rRaVHuIoImxCoY9v6sijdzPE61hXCobDwhYq/wJSx/SyGtyNTdkyZNUNhEmtgyznK79Il2fcGcY
XjSVTGOh+yA9koL1GXX+ZTxtBsZ6f1ihmB5yRgYfv7EGTnyX8ehP94/H507OB1B0LPuckrIhrqex
jJwLd/HoMcnpvXWQeI0QJIsJT0b8Kh80apoXI3xdgd5ebFEyjBxVst6H0Lx7jgWh4kt9IKq6tvDE
7l0S2Fxwr5Cx5TyWOkr7QqT6yqxLGVgAaFLU6LUuBeBBu2WMwB8a2rQuPc95xbFQUIJOaFSDKap7
YanbXbfy4Ip0xTbshkhlOGt6VqqZEOu539XgvAWrwKyLlXEo3CpALPDjX+G1jdMA0EDcxSpPvuFT
WGArirxSoiKvKeY4aY0urgFcGNnjurHwGd7XizM0mNs0RIkx8Mv5fiVfLthxgC8npI/CVHpL46qH
HrVKxZoEXumm6l0ch3W8ZA5Qch2NC2JYHTEyNE+7LG4bArAJjEZF9atE0S7jPsMdvC6/NZ/fHghf
qgcUuz8prQW54voCKzuRQ0a/JumvbycNk7SNevLJdomNRPSiZKaX3i2TQ34MZptuoJwPJiVZ9FEy
5tXRw/xUKj1Mh53sRPX6lHXP866eP+2W7oTWVAhX6FIcjEfgOEfeLG+FUO8AXgyLaj6fg5EFcE8K
zYx6BOxZOe4qDt4ml6PMdo38zQUZgZAHAfCaJw+2kM2B5usRblwxkZV0/zJ1qnvwACsj7k7tUTcs
p7Pc55mXaq4rAMAGr6bgrnEzZWXXaqVZDtmcJ3lGgksYmLISxVaGFRh0BS7Pfk357zeGtg6klrCV
Uj7BSlMAwZ7r+6WZzCtuToyEJsk6tCXqfddb7fa3DfEwYzRPBk+DCnBojFf7/KwfJRx//x3RTa14
q2H6mem2Yg505YCfrrsHuffm+zghZYDU4ot0340j2ptMi55AZM1omhgEENIwqYcpEHkGRc7ZxGsw
1NgFWXjzLvpxhHGJzDDSHyAbezS/ksM2dYUSslLnt0mN/g9wU0S6IzPzZVsFecQWSTBdVHZdqLUl
Khb1htTR14SdNun1h/tQSH1Gs13Ja8UEFKKB2kjM5j5gawoxEZB6GMfbNiPqKJxMoIe2wvI+7epd
u3yqVV2AQwVp41YXu0vvWNHA97LcogyG0hkwRxnerfcWV/4vIMsdI82qd8DoGGfhz0OtkCurlkR4
vuZ3/3k7VfuxohWFRy/crskjW0m0WMzm89sPHo7Rulx6UmNtS0G4tg+XvVG4SZAdM0UySdBcTyPk
0IZn9KrVv+Uz4NUBM/9O7AZPEIQ3EkEFx7Oy7jhr9FMa1V4xhuBLMWRYjDnZC7L86ejKqso+DB7N
JnHQfnBZr6FW6TAso8hZh6eKlYBKp9RmlSfwy/6VnjGkOSS5us+0L3z0ELmU+5r4fIwmRqL6fJW1
1EcmgtHMXP4R5dgYo8QAF1keB9fW1ax477xqrN84kj61OxfELXUM9LocXTmfuKxRX6uZEVy4UZ5C
00XJf9nRms6SH2htJ+myJ5hbUGLmcsy4BSAkZiUmUrU6ME5YWaAt3brSGJoiuA9IVF+OJlL8WY0C
S3dTFs0zwZdtJjocZkxH4oNnsnPWfeNFvCiJ9+Zuu1owqjb5udxt8SiE938Qbt7leMmdH6aVnBrb
Sl3MD+aaHBbGbc/ut8iO1uD1w/ENVBqUUjGVu/y9dPWQW1Oy0UfSSgtyZYiQgaK2fwLaXD7cyLOM
PZnQXDNec/EUm7Adq9nPiVeF74gQ++kgr5UQx4buBoymMQnCpmJQL42yQpNe145U+J3E8ux+0ymw
HLV8AukaG93aPeWuXaeOEMuA7ZCeL+9hcqvWmj8vv6berS6bmO5Of5CtzEYBJsj9oxLSvWmvP6c2
eQ2yY3BebjRGExoRKE6Q31nDljrSn1Kve4nNP17DoG9JyIhYvzqe/gm2o46xv3yk2mxSkRlfflc1
vmzCZvEUTswZntob2xbB/moaIiLfwSyBt72D5rQ+o3oAeCghR5xf4YriKX0UY6enISZdfz/gm9Zi
1nmDOQ/aHr/xVMgrW2rIB9yOc+O3dY1qK74Aqf/wMpt+22GXTdRO323LwK1nsU8j4ltNsH05E5Bu
RGxm8PudkZiwUotEAUZa1tx79zbrhMa4aeBMFiMsA8UR7JbXV6bsiIaLzxc5q8ZA1ut9EA1Rs67H
tPzmR5K6sQLzbIBi6o16lYqPSyWdV/m6BRvhRE0D81Yjlipw+PJvJezowIwi/x0c6s7spS6usHgD
LK/9e5SOgJK7BzZK9m57zyEKstazBo2GuMShE2WG0OKUj6jJXJey8GqQ0spc333eAoZOuk1+uwXY
x5VtwhKzbIqaGbNiE7+2O2+3WuGIGtEWMAnakAmoguYUURSKcnz7KAVAJ+CDusRqO7mb9medDnow
mickRJTuxayUE8X2JhftPMeSmQmZD1tz2AFElZw0LIHxE9P4rOXpm2fF9k1f8S3vuWej3hQ2fgxv
eRQdu0LWyT/mhd+pGwILLmdsCHvB6oC4w1Mzv/woiyhIpm1rH++ljbo7S1bZmOl2Ull+WfVyKF+g
YxRxPX/RmFuW2Ha6Tw8r/V19GhDSf3kWk7l6QmWO55urbHVUeZiN/Vl+WpoO/bgy3mkUjuQIIQJj
yPjMe0Z974AtYrODKyLDnQYp3Z2jI/W63keKanPBRENBZfT34lzhYhoW+zy/zrYrCGBTc8dV7HBn
l6xJBYQveGtTLh8YcUcqaBEPpPTkR3Lve2z9APuJahCLkr98TpVQNCAAyxqc8ZCQJX5nCtL98guK
XXnOmz2IyiIHZB6LgCfbAqhbw8aUNubFoWejIuILFrFvErgMZb/PP9Wy9hN9peHRXiN50MoL0pxz
ciwNJsPMDb8l/TljzynJM89OWDlvvLZfBWXkydYD4x1gjkR17tIg8D2s6KU8Whfy/E36ytuBdCDH
3BamvVhFvfG8pGa+IGXdfO+mmQCbJNtwsXVxB8pZhJSAfpzHZ282OCFd9acmw9guuC34s3F+Q/Mm
pvqrThzpR7AxNW/eeqoAnta1CF/GdphO8kh66JCuVNsubHNHAR2mn1Bpwr3vKDvIZEaq53NRPIq5
0sNMCVE6q2P3I4PqFtIo06ycxW4+7xuswG8tz2R1QRva/lUWIZ9LnmdoZJlM8zFWts7aJQPIFQmn
wDARQI7fiXTy2JNYGsYF8LGcNAgRHPaBVILWNPv3cGPFn6yVwnY8bcIJrAh3LTuLm82vR56ouc9a
jOrIko//hYjUsxkIEgk61LQTW2pNOV/aAgmCbuX7zXAbRxoubB+SW4Ch7e5wsoCI46Ag7TuWU1rc
Tcl028PM78Rjf2lMSX+IbNsPpYWXzncMjZwd9ir84iR+90dvQAxaMsoQf76Dw5Cst0kgM/FBpA0d
/TP0b7UfcSUZi1sUq04bpFLSs5X4FMA9lvXl6kazKUtdxZIhKFA++ugs2JBcIxumBJqfxUL1Ce+T
ZYPBuw/qkId+cTHYIa9lj8mHQo8ZuHUuQVkSiHEy4nNJ5KHXXrhSWAaAEPAaRaCy8HcNmA2onAZi
a2lKrDnL+kMSU+kX2s7xUCaIgcqSbkjU25dX2k8bxAehDL6XDpBh/f0DKBlq+ip3gMPfveLTn1kx
y2oMUH1DZLBZR+ojv7GREXRyB1MhUlKTxTHs93ms9Ilc5VprFvI6oqRUpGCQ43URxUlU7/23a5OQ
68koxHvmTvISGkWwkmPq/V0G9C19oZRZsspJ62UG/MBWs9259f5IXt72LJw8YwyyUbJh7mHQ154m
ErPfji/xeOkoWcEGR8Xj/5bOmBaxxxWWhq8CVapL58kkVnPPO6G4GkeZOUOJfEoHbFLT/2wPYVjB
KrZwWUxVp23btyR8vyurD693TD1gOxNCMC5y63WBnTeCjlFYXEXGRSb0iUflUvw4m9M9MtEoSEll
CAk/XBfef64Aph6be7QUcAl8uiGS9iYGfCvequN/+re3U3PDWGLwTwS883HgFGpVFSBcJEVZzYGb
Xu07TWk9qhA3rlhD9xs5cIP238u19neabOpTz+c0p0enQ8oLxNZuLeyBHgFRTogdER1JJ7LA06Uh
/JsJO/eMNX4oAplPnh0o7KB9WNll829E4rIV6S9jzCyrAX1reErjBtyQy38CQzVsz6Tp/bFQ9VlP
JIx4mpiJdD9/s8rBGK0e+aj0glh43NjEe3eCgiMI1N8yBWd/HWnQ0Ltl44YEwU79QP+T9tuJVGAW
CYxnRUA24yTGwoycWad/f9YB8VPU4/w2ggS3/LgReCOziSIqTmyc1vU1JvVtT1nLC3hSHXR32rOg
5wHtSLTujW8dK6oF0PfeL2IGKlvVpjE1YZ03dFRFP9ObZag/3UCXi8PTja5mFFQPR6ujpZ3j42DF
Hi/TUK9xV7s7+CTMzpiTtpdBRbXwADQaj3FRFZyrwXfonQrOd/7izWsXScW4URso2p7NCuptR2n8
9V5JH+Rxz96enLfc/sTAgJ/eVf5h9MHQp4bYtEC4LlkDYKauJZlS9KEfGH9utnhqCKSWumhDPgxa
6nCoS1l3+rzTF/JMRTc/A75BUZwFUB5Lb4osc/+wpWOLlLYn8hR59Pk7RBeWh6odendb15wqCyp3
NSQspox/tWMuxjGedkkmei/j6KGliOeLT3aR70cQds0L3QQCej14gBg1617GhP2TeoXDm8k8/eOD
E1Fg0k1Vr8vzy4tHW2X4NSGu7ADSoGEFRD72ySQrOxzPHP6FRNKJy+dlq22X7e8K79YxT7dRZxA+
oMCrRQibx/wKP1PqPulQLCUEJg0legr+bg1B1Ko4aAJXyyvb59cVexTbj+ztdBY82EmJ5T9sijPO
peW0DMRIQHmLeMpLI7E0fZaMACId2HIHCbnb80OZyR0xaQ5RVVGfJ/hwoQ31VtnIha2rOyTo/u2J
wRLO+SeFDWrw7swA6AKONiElEECvGD0UXBUhInGVLOGIqJoUidb0LOtmWoNET8spCW+eFfN26Adq
v0bELpBmxOmkQ5il6SaQTbOTMRqIzwGTMrxHzo+PRhICvMEwW+MlgkJbNnKStDV8Rid2eUrdbHap
cA16hHrw30IyaFaiM6Pyq4rrfnEWOFX85nDcwHYys+Ny8XkqJzYH3r+EwrpDOpn96/Fuai06KrWz
SHZUgD2tsFKjzymLrg0jwo2ERUl1bpPuPLRix4avmsLHazc8G3UlZCAJny9yugFyPITdPFA/vtmY
9ZCEyJ0i2UyAYTwLgscH3MYditNJRHAf3CvEtGv/CMINDUnxGPvRfH/YkO0tFIp6J1X3EWsJZF7Y
jn8e2pskZJE6JLNGa3vUow3rfeECEmmyVnx7BCQMsrEsJhcYCtUjElcgq7UGZkaXxxGjRQ/cQutU
o0ob2AoDHeo4L4EmZc8hi4Kaj9nme3QHlhegcNKoLyfCc7Dr2TEX9qJGPw+g69HiS83dk8Lx6hXV
o5iE7t/MajMqrefmEhJbS1izy5Sic7KkoJN9oqSS4Z/jIAgk6HqVp7AKBVNf2pQeS9lafSAarx/q
U9FkSWI04kj9snPuC9cqb49+fDe51xHbt74GLfVeuneGht+dLKoU8s1Y1GUwzb4QsYkU/6mUdGKZ
UCIkEx1ppKpX9WDbkGu8yb+ndX6BUw79Oc5WPaKnbnDGDmKuFZGAvCI+2AOBpdgg8GFLNTTJcnN/
Rt5VrwfOIryqLHnxpDqesxCmYfu/m36U5qbTt5KDybeNQYDvdBQDPuj8hUU7prgrUmrV5SFfRK3y
rImI79/Xr2lRYL7qSIgvc+MWMcxihxlZqUk5td8fEc1SlRHJStr8PJXmIRDlM6Xg9WoNFSlS2niv
yMsLL34OTmhD/lFWeQ9nT5N/IX2bYzl+69CAU+DxpkQM5nbOTs2cVO/2KUCHxLVlvl5IPE9OrRqw
ncx34IwY9cCCgGLnmmQWFC4dQhA5YJBb76LIuFQDbI8gH8dN5oWIFaQhonZAQPsfWdWqWc9iRcpn
upo1YUp8ajrBXBCda3A5zR1frTmZAvpi6IfUZeAh7CPOMECmLObRbuMh9uhHI4Qr1O8yJlUaFHeF
lpPt93tpJrX3++6mv1SlOdYnyHjwOaITYWP7IgIR/qnLEujHugqnnC20eYevOTuXozIBSHpCZw8r
iyxm4Ral5eZSUtq7JMZ+juvD1HAkbOJCXzmMpShJxAl6eK1W7aem2gShRkAOhnjV4rpSqs5FLIkt
7iV6z7zv/JU33/Ysh9LRLqJcixI1+vlc+bUQADgYSkxy2og0C7j0NBiRCtgoEEe6dg+ddZeN2GJy
tH7tl/qYQ+zgrBS4lQ9FlmsKlYJZT9TGB8INLf3fZlihL03mdhC6oWwFssY51J1pZ+nKfTvMH70i
9/NkXXedU8SKlh5nJ7MMSQTPTBv3+MEj/iHjxFvvEbsrqcf+4ujeOuRd2PGzDEAdtvPN+dNRUCk+
//xuBjD8OUjW/goRJqRGAcE6OUMvufzeR8/uRYcRC0UL9mo4aC6gXi/Js+aoDImuguNkaxMWSRQS
m/JAlYWR3ZqgXEaOXS5Bad7ZSnQoDQVgL2bb+6adEm+jLm68oxthzowiDEuXRuGgdxn/LwTpYC6t
p9AhAESiFvJG6vhFImNjrQennBrhUt5O1uJvlIAdDPx01Cw+NCzoq8Uu97FauKG10LU/pefkVck6
Gl0BuhjC/EpYX3XOxkB1iK0suSwOlGW+4mZhS6df4w1pDal1ZYYMYrKidCkT599vuhm4ANimHqEb
UAgJlWy1eYyLlCZhCk8PQK2lRrPCfJ5NzcC6mGkvpsA7lHzF0T1LunuE1x6/AZ8jk66VhMH3OH5C
aTdFGXTedc5cQYVzdsDFuQ/mgO1wBnhcYbdwrlF9De1rXSruj+CNcq5ewV5etwlKEAbMHscLDBQ4
BH18I2tDpwvbXWZP1Gp7QQq5ZdYj45HenbFxqiz30ch+JatBQaL3JI2xkTDyhaF3HIT16q8PqkXj
CAdinrqLwKHqZhskkbNH+o/cJMHWDYmwVxH+8yD2kl+H4GLff3t/mUMejhjLse6IdJgb4jrhlm91
pGAdrxWd61EshWxoJWgdDcH9MJJbbFgwlhPEWeLRuidNeOMwmysSCg0Jn/9zsHHb8jLa9KYfIvZ/
V/zmxPkTm2TI6VaoJkEpMmdBwVofRboPQW6dcLuX++Zyse6B0LH0Kt+oqrH0XYAkTv1xiM8Osih9
N2LYtZ5QZCgx4W6b8x29tOxybq0mmsOm4IskCsuC7Tqs1jdDd5wuKjy0dMUVNqD13EJzys0sor9/
LY+6qv0Kct2+/BCgNYiAnVk4Uuafayg7gQSHRkug3zcrB4VMWtELY1I8Tby799DWAXMXgU+XggbF
Qk6Zax0ZChktcZLQfeNYsWufEZvvyMJavp2PeNg9EREJ09l/kIoVE6/feFY1L4eaXIkF+rO4+B6u
dfbo7Fi00tSqlM+ECeala6NmkQ3YCJRvUOZJQjIyiS0L0Ms1jha1VP4EYoFr4bEdolQdwEkMg/LT
/hPLhFvKemC+vPaa2D3rGc8w9IVVxl6OwgzHS5ZCMvNbBGElllII9IiNnjx+ZZPhbn0c4RWLixkg
hhfGDet022GCAssVwj2R8x6Y+DLbxbrG3Z7usXgYrzuvfuRrz1odbSY+J+lqfe520mf5+wYuEdpA
agkNmm4tkddy7f3hiQSH7rbRRaNBMt9HOldGrDMFXcFlXtL+6lbGFKy8F3xHpPF834kyt9ugP42Z
BnQFZnAUUepIzusWdIOKyXLu0UI04xyciifmWXky5ZTtxbwfDtW/uz3L0qIrsjQhYRsOuP9ODgfC
qfva6hZmPCwHUsX2cE68otAEqz+H/7gCQfHTuX0/uVtwHzKJUUwyxgHLcFQZdzpRjXQsXn18MYcu
x+fBPCdM74kyMy+OeUtTH6xAB7NO4azNh4UINs0tPUyI5zIlPikfCBxkjmJx47CulIo2xnyugDyG
MzHfZPAn3jUFdCxh2oVRHXtlk+dBJwaJHmfYy2pk7UeuhA02O549aTGPT6j8q5POcK19P2FtMYLi
T+jWMCMo38kJ4xNAq1TPZmngjy2aBaCMQREzVtBgaQ9WuO9b15hhuolWDwh5egJfwXWrz/0dgf5L
PdpSYI3HythwLrcDU9Clfr6yW/i1BV9gLsUU4FI4mQALmQyvqVsNn7lyD1dJD/dX+IUNE8X22xkg
HKQOTIENAtE8WeIwqeUDk0vrC3r8F5T/BKtZ3AAp21WgjVbDj3gS5r8rYW5RCrKDYl87FSygn2Wr
gt8CXUxmDgMd16rimb106R9PRMfbIUS8ATKw0GVpJZzneu9bZy05UGWVb9g0sCwUxYYHSVpANWQk
MXB4woMznxY9vozuRKktxaIRRnlyCPVQ7V31Bdpnz8lp4nnoq+SSOmnYyjTrHlW8nJMOLB8QvHOW
xbHuhFbWmoDobvXXW4+PeQFMT3wwf8T1jnwxv1vdYnYy+LttOyHnGw9LBTJbmPWTTXTMn8Tr8Mgj
aM/PUMcM7QfWL2XVlP8Lygpx5rnoxF9Ki9cyBtoDbt5GEnR/2PjTdNw5m6sXIXLhmExJzCoZu1xU
o8xoMmtxwI8/C0dDG8GztBRS0phRFTbMgms9jxUnQH60MlFjVK5LqXJ5pWzCiEgt0Xl0YA1QL8tM
Ez0vUq3hYIVUE9Igwnlqb72ANPGIXN/IsvNh4KpCm67+8FAhQgTpBKmewPS7pCx1Pkl8wuQtAob0
vl3TmTRN0+d8H1vOfitNI5QlUw8GQwaOfe0xVeW4wrqDQ/Z2a+/3es/RqVvbM2Zx5Ikrk4hUVZMr
HgSrnhhjJyfHuWQ7BZ29fRTIyaG9CbeBAHgRrD1lLhFOHhUGm7UqoqhtwFCFV6WQoqYItW0jL3eR
+vARuWBsMJ2wAvvWf0sXop500yJcSVy0GeLpqgawqKHirVithsVOxYWqRH7bpy5mjd65vliT5cUB
AsCxgGqWYIKfrow+cj1wBBLgLq0SjtRjHPOjjiL8dH6ZYJXI6zTTN3aUjOLL4bWLst+rkWrfeuFK
b5JjB+F9tmpEUrBdRcy30reQz3qWwf3IhXppsugDqB41iJmzDpk3i3E8uxuPwOa18sjdz3Jvk8WR
ik7tYAmFi5kD5+D17gqaWeIi2EjlUXM1YNLhk/Pw2xDoIkywOpj8pl047zJ3GSguZv6TyfOhNPkO
Rd2QUzaKwtdj+nkcC6jHaqKqqbCOUvI6vLnAiiYId9PlQDQVqMWGRXEtA7UY2w9oUsOlvDQfhW7Z
OjwtqbvwBmN2HuW2BbCnfIyRvygcH4NLYW/kXeSVViFWkwJ6a4e6y0CwTSP4qp3Ol4wtriIF+HyA
K/dg2focArDcz1MRJsv1CD04aVv7YE5H86+UsdswLFyCTdSq9AqxbieLKWQLEMIu0as1rEqIklul
HK6nXjv/cKtyxO5AdARaYfu26Iwbw/dEexm1z7t7q+8IxQ0aTdm1cOu8c4qF/u9jI6CV3I/lzyOo
nFvRLygurkH7/AFE16SHf/pf9cCMxprF6RJ8nqWGDRW3yO7rShM/pjrvsEleYIaGRCgVxA+JAFce
zk5ZqkPdZfiiKSMOrjfa2REuGN2IGD5F1QhDnKE/kGGo6ZaGgtPDlFzEnhE6Y7LR6wVPQZJRdQmz
pU/uQjy5EAAbZRxwP1PN2cBfxqO5yKCt19bMJe388YMsyH0JPAiyheifVSeLW8zH2PJbPcwUbGSB
6d6R3azGpyvVIt9xReS156yiuNY+t1vu+WfZnRTnG9KjqBeufs+rGLOoL1J37ItJxqHNNUfCMS0b
/Bq76xh6nVh4OAZ2SzDM7GOPrJcwsMwmfPGZ+RZzORrMbkaIFqHYSa2GGqXb2ZFd4RKddjZtSwhN
kxBoTW4hvp2+0U4h59XkIbPq1RWg3bIdLwNv0yOhpD5JWb6rbjDODyT1/d2KTLfWH2ERGZx68NG1
J3nK4AfgzLa+I5zw8RABYWTd1myDIf2ie+07hXa8I5D6gQvw6wNcrYn9nF/CiclPQDZW/vbsFt+D
tm+ijEQpnwlTuDW6ENeb5PlN2o8ksWQ3srpG0XME7Kuopwr7yUt/wuy4CdkcM7NHWvqQbS86ece3
3fJQJVyGuPSr12s/L0yMkaIagnZ/1u2gqCaeE9l7u60wgFz1xIkvhrl9Dx9xYQOD58qpfBbYWEP1
SvxLFGCuSh1wz/86SNWr8OjqsXPgHTG6Gfzmvsuv9L+2JOzXFZI38VyrB+d6H+xHFP/o9dQIHUZK
JoSm/433Nr6cUvA5MpTS9d0zoWtwXvPtg700QimPEydvbE1ttnQUnFH7Z3+8XF5t+m3m3GUSDLEe
zvB3cVdP+SyFKSNHnd23Odf6ppDMHAeVWYUmqxoF7Xze5joN+qgyw8QDAt/NPISLBRTXpAGlmmZn
tTzKSWfgAEpkIkTZ+AORyji8o9pQ6mEKqUw5EkN1EWdIik/pTNuNQmajN4LkHrqPfrKFJt33cvPi
APWUH/1yMv64RuO+7SlG3w7j3JXsFufUs3JyiiId/qOUXXEXlDgnfWgGwBUWPnYYfaSwmca+Uoep
V0wDYEf2HowPxDfsVWEFoq7vTqBfT1jTSmXnHdcJjhgj4Ham6cJdGi73vDxzzcl1pKrZdIHAOtVo
rllO5FQLORazWQsO+QovPVadxlrCryXtEa1QO4hMIVYue4OQP2jLRVQIFcehC5bdE2idX21g+AaW
6HT5VN2rQWyt9IdsWZiLDY1xGYG/dYtI5wfeaqqnVIdU8CL2WEMFhdC61RNvjfbVdlHAltAWIVVQ
vWdmKcRbOJ7w4+8mzqIMG0LZwVClXCmsKDvZOHhQ86z2iq6cTzBLlEWUIZFpYx2TnHTKumalLxLV
awaiLtJ7JHO5X5ybSaKzv5mOpE+MkjkKwU62WWHjO56evpB3pyGRb7d1/5bRLlK3nb1z6FtePOjv
hpViBTdGizZiMObiG/A6yw0H4ZT7mGPcpFzs056T3WfDP5DegPuUSiY3j+/ivH4hO3Xx5iRz+Wug
DPcXyIM81MY1oxbp1ixSWILBUOz4+nrjTSPtvOuIJ6j54V8lruNmdKJAiMHbWD4vuN35jiuhAHCx
61+tk9Rg38Px17BN1cXKQbwJ+ZGtbhxFobg/GXisYCXwD+7HfEYFUo5WHBerqcnHbym+yQt2SK/d
g3+/evz7jXK8aBeQbRkw6rJyL2Z8/qxM8MuCkBYAD959n9KsBPtNs83dx5Oeo/X5bAsNV8LBkdfs
I926xsqWZEgjqJIo3YlAXxTlPVyZ3su4nLKyO1CVLq1cSWDZQ5f4CJIq85MOs0y3tgH5f+ZmmK2w
poRJnMFV+pf8nBQqEMrh/banoLb6ad20Drd7F1yJEogyKF/HyNzGHhrynFwd6EhmBN718aLTGgBs
91QTC8pgwySLDSMfOAocKBagHtiInv1gSz4SDYmtbsOXMgQDvHTaIKdKiqMbd/YK59Mkov9qFDgK
/kmvpY6nrxKcdnxhs5uGnRHOYVCZ+y4nflZS+370SMfsMvmk+Nb9ieLYIC5vShybfS6EPbM5Vr24
8M/27sNnGAOLE8g6oYWLp3UEAWhImsAuzvNOVvhN1EcjmgR+e1tzEgtU/l2rHPJO7hDoAO4ijoEk
vuTvNN3/907NEyWAFqxOJDwpMpFoAM2MhfLHTzgpkaK8QqTLJ9owya4l8PPOddwetWjOwpClScnL
mb7X8O8BD4M0y7bK2Rs6hke+PWwN6yAaNfLsxJONY6ka5mmDpDANLYFj5CamuHs3WpqV6s61yETv
jg4hav2MjoEJACIl5oy0X6IyATdR/sSPD6f9+IfORHnwLLp8kRPLzusabRw6yQGXVKTJgWcOt9D8
giUFdUpYbYoUs8k6Y5anprWeAErdKf/r1lhQ+9De8frcAGSL56uF2Gjw80Bcff7/Vg29ZOeMlcru
r5OUJm2Dtxei1EBl07GmXz0JPMyQtV0nzhYuO6cC3eVbg0xL02Tl9H9FoH242+lSu4X4/HRVI6pA
rJNVZ0GrQBpSgTrjFuT0pwqTWDX2Ue2osSeOjAHL8u1YkD5ijeEBVLNdyju2UVxvOkFYh9SaBkvd
0Ga5RtbFHRRt+VY1ew+cvaUYMC6gyvc3bGy1r74csh3vY66ovBOMLQaPuUk3FngjlestjyVgHIyf
xB4EVQ75UIMN/kdgDQ2t8XlnXJPg40qKZKqreOQmQyPyhh0xl7EHh7bPA5vGnxEspd6OQ1TO++ME
GN1KOVZyinCcqlWBBtx2OiUHTDO8aI8TZuhkt38g97i2ZIizx+gFIiwGWsk2NdWb7nJGiMUHnjXK
SoDAX6v3dNMaeglXjVA6X+PjwurqqcAwr2EfRFJdAUNbptRrQL0zwdufmd7oWhQKL6K+SGCTjSW6
W9GUy7JLfQFjh6S1qt8lvLCL+T8YeVqcUYBEhTqgwwf1fYq/PjLeOadrpz26sA9IL0JjMKymiC8/
ixEpcoKpdtwadOSTNf/rZuPJPWRy7zabXol5/trvWC3KiKrN6g/HUPfAtPodNXAD6e3FLJs5I6mq
s+5/q0wtDFr9CCz2rKbvGQfK/7Gvx75JIWKFUxd3W3/UNp1bNxsWbYAsoEFMBugO2GeitxGIPGSO
fJuaTSCaHKI18zorEX82/8C/2meVFJ+akg8n29lNKE9P7hiIrvNmVh4oWQWynHxJ9WcmbH0HBjzx
Yh4t43l3IJTp1roPSAfhGlBCN0g6fXtvVbhe9AFbjd1TfEk22nEB0pwuVJ9soFOeFjNOKCmZ+VCn
yHoBzdBJxfvVnjYep8DexvVovCdUxWYN9Wf05aoDUMx885IySyOlaWn6hNZ5yzdmPyjAIinZyQg+
qwzIH5jhd5IxKvsokXIroCfbqGV5ZEJPtG1s9pwVPjtxhn7+9Gs8DeftExkzf2zfurlurzPy+2Hx
TbC0UuX3Rwus7gkSRRDS2+Kru30D3+kCcHpnhTORhBQvzEaaxhoixnT/NlaFysvf3Qo1gSrtbWML
Gp54Dm92n4InyawlNFBQdfhzbdqM4wiq3p0YLAudsuT7wNMhIfSsO6/SpKEYKbWD3WDwDnn8zecc
QnWExh/i6x5PGYsFDHVBmwo0T1P3T8X+c2oaFKC4Xc1KcrXbgVGZkfIXFwG17bfiNt+ZhUAdBSms
DbAeLvhh9PrqKNC2ZSJRWrZV5v7isquiyOTP6OmDJ/QWRlDXfOqkOxYzV7V9svcx8mTOEuiO7vmw
jg7/fJMplkvOb2SGMcyUfeqPf4b+1LBiI5qpyWvzQiQrkRbATewaBUDqQGgpm0NpytZykHdw1PcR
Wvsj3/v9T1bsrJUHTVm4dbVJhmGG7AKugEICS5UVhKXL/lFMkQasrskf7fkuUPEW6Mi64GazHkV9
BsY22h/lkEI2+wVgmujp+Gqx1qGR/CW0cwe5B3kX7s1H2cSapbuRwDJitsv1fFDr52nbSzKzBw3Q
PKdeGZQBE0tTpWVPKxUu9DeOUAqEZ3DSA115bgBW00yNZLDxfITNxkx9pnN6GE8+0MMDnlVTS2kF
R2AM18NLZLJUrIjQorpJio9wqqHR+ZKE0PK2+NIKQOVsXDErTCL8/BYEIdYJnCxYvP/Idj3pcSAA
hTuLSYrH3cpr8IYLffH6T2aYVM2cCrCR85TqGn5r1qgw8IsMixLc0p0T7Fdw/TJkStdXDnR+78Sw
cSETjtAHd4m3Gh36uMmZIuTSSoTrSls1XQfXbZSqpQAnhbvxY4HCFOLmwFTo+p/c1pyuUadQyxIS
AJrA29rPV3MWhdzHDdclQsPE0Chx90H8Q4qH4Z9R7L7FdVdW7cDZ724XSH8iSfvmoTFx3s7p1iN6
IMgRwECu8Y+fPAy4vFLu5squoxyWt96eK5Zdbm4RpYOUrsELhC2HK/S6Fvx0x79+YYQjsWa66sL3
8A8Q0e7rHe/axJ5x+JXrrQ/PaloMqIO9VI37SUWWpgKMu4f8fWFHxW71V3qH2+YxomrYic/YmxRy
10FTzMFW8+jgc5s/jpFdY8JII+uXmaXLKB9r6Ceup1QYicxaFhkSfYByRH1HCu+zMzXq2U27sMEp
1yw6fIp5NqTFeKZpK9Vd9OAIlXAynZoeCC6pLBQKEKPeQv+Ebny/iYUH2SlqzAcElJOmMhdxtnn6
OtNs+zeEMI/KbFRPt5s32+sfC1aTGDW4ekJsqVJj8rW4uw9MZcEg/D5+w+gsv04in/5rMz3M+cz9
nHmpJTTrevxIDagL6Vn9yH4Vb1wKTCZh1/rthTNnpejPvXhdIefBkC6cFC3C1PorHuh6IvMm9RMQ
DDKMscJtmjBvPCWULwHHLcKxRA5KYYZGmbPbPv+mS4k5l3DasWNBDTqfjm05eookSQVD0Mc4A6oV
M3IVepmrEuHuM3qrT7V3TqNfdlGwjNmSvrljb35M6oq2WeLwzI4cIVCD5tNeCy7jY2Dzhc30xKfD
6P/Yhrz3grxCgtjV6wt4CTFamQRidgyjCJ14HkH0WFkCjwvlrlm07dq7tp2pddsjF5Asz8zEUuD/
h/pXqy7KLJuoj47YmFUfZTZRDzjFRWhoS9BsJorn+fHfu01UXiGsbBqeYovWshgoovKaxBBzyIDE
Qjga5je5JZwA5e3li5koihncodMOncR3qHcQcNhM/MyGB++jNVeXFBsSo3i0t0njLS6XFCqJv/Ex
4Z9qMnDUW4SO055gZZM+OSvwsilWXTr7DDoUTMD+5yzs6IB62PuQ5lklaOxXHY7V5K/mOKSKWlFm
bN+J8FJZHAmR6Q8sgNs6Y8aVJNp8oQNN9dE1LZuLtMiy7JjzRTEl2HMy04s6Y58JENqOcrieKMkS
foluvB3y/xBSVBI3O8kyCtak/jAGMGhQsJo9KZBc0O1xz2Od/4arenO9oVm/J01V1qhkZSO0TPVk
6RVzPxbGNJ+4ZkV7M7M+Xjri8A4UbRV6LzrVBcyjYrlromP4U+/Ravnu8wzFDFXUr/SCrkSWr1zv
BBCVum5co71e5zWQQXhbq4APlOnTNRguBx3Q2l6jYD4uPODvzgn5L684unvoBE0wVbFq1DGFgNS7
+MDYOTxEJyroclEVJo4jRkJ1ezRu+y5iDEeQtPkMX+Eq6EK+0CKj7rll4IXmmv4xIJcTDeBjTBBp
2Own2kEbweow955ZcB3uVaTdpNVyD8ArH5xNejmU38vwDZWp3/Qwtaxipugx6fBycCaqL9lLD9GE
JMVlRk32694cHxFpXK3kEEqrjqnbZ/SJgrI+rpKVYTCwGbqjIjA040qSdufmHhdild0EZB+Wn3If
JIS+KguFsLgftXlUOrBBBaJfpHn3WDgFkrAi9znxRKuNHwvRiqvPrD3oRDURFneA0dH3uMl19mVg
RcCFbDPgXpxS9QTaIwJjJ5DAnd8RHT92/5ow65toUmf7peJ+XG1aMSA6j/HJwBsdHFy9avAG5U4r
RmVmvq3DGrozQixgTpcl3EoFTT3WxzAL9iTeOAw5Xtvn8jfGXD5igj6/3IG/YrOnD6oxAE0gjb+s
npH/OnR1+/1cQQYP9SQsA+OVfC49mnBA0ybjIw7rtHkgwFFz/mTCN44dun9ej6VIVgIhBBHWIxc8
NDp6i2APGqwyCpw3WgmZH22xcVjR9iLOVtSH5IGoAUFwAqv0/DYxGVz24/pRGbyYbgolDHipejIg
ogJg09xu9hkbhQKhFegUVvJ3f6w/KhIhXVJHkEOaiI+ya13sUWNueZBMtQtgNMr2GuogL7JoeBjn
HDBytCCI13pNZyrt3WyKU5a8iWUVIfOzJ6/yNET8W1yydk5qJqYqu8VhZVgq4+61aCcoaiRKKfVD
PZy4c0cFif3esX7n7YoDWJVXgkNbTxNcb5YVt9pW7bpMXIo41kbWgpfFVSHOSCoftGPIsWqzmHDC
WADF0KZZj8Kv0/B97/tV5iPN4+8tOb//44uRwFdP9F0Cl/4HCeR7NGOxFsav03yNZPVRBnESUzxq
ykPz1KO6HEViT4/QcBew3lKpGXRIeecDMogptfNtmWPhqLj+VtLrCTI6CNTyxwPZZ1i5EAa5dB/l
ztaox3M5R69ICnqX5qGUdJnfQD5cTP5QRWrkPmhz3Mp8uEawzeEvQfCwwhYbHc2gMKeqSKXeIvk3
KQLPeD0uCoB6E1KSS6f1DtoT4LVyetCEjlf3rqq4wi6vzq126WG/P0HVk+W0ENfQvTN8M4VQrIoF
xzHPFlDaxTEsUyD0xgNAGbWI7o73M4AHksOQ4jmjMjko5E7x1epmUKwH4pBXaQ6UU3IYbgmsvHF3
+2cDW0s0EOe+VDAvDB7gMHskj3OgV+WUdiTEtixPyZSVGeTlF5+xgmvT2xpQnskhUjrdca2DlurH
URnIj38ZQ+DM9yurPsGuy3uIblLiUt/v/v+nVT0A/M1GfUyyw26NNm6BtzidQs4uhG8brkXCePBJ
3/WbKVJGzn7glqAdPb++yuAuj4IhqTUpJUifhMnMQb/N0HW9aPwJ9Q5aCf4lvheuJRg17ySg+1Ne
8il1iZwOwqH2BtuIVTx96Zh6Y3FMF7grxTtsrbkf5D7okbDDmhnB+2UJhFCfgW7ByndIbEAr/DPq
WMQILQUh/bl+Fnr0l4cVzdhgKG77gAVVRvN7jxtvcCcj1uGhTkPZsX+1HmnsvF+aO6AHTyK2Pdae
1pPterS/Nx1eoiiYjAz5IyPK2WIfv4uIsdHTpwMwAEX+xgPtYA+ioPt3naaebvTDBLwjlz02f25Y
ozs7rMnueVL8F5rO9/LpNymZabP7iBoZKpsDNFf2k/Ug/rpy6qrNeLoXBjfCXThs/FLgvPff6Da5
4KybEuJXdAUPtyDz5luap2SJURTyEI7kagnbcbAaOlHb/8iGRCSogmgDkk45EcdDBr8aX8S2f4/a
teDDeyTUV7B51czX2+9PXKb9CfaRNQWtXf1fjPkxb0aROG78l0NFP4TohXANg7L6LZCkTXs2G6Ex
9rlFnEE9HCJkegDJe8bjsS+qQ3DDpV+uoEUmHCe9TEeXcv2KZ+qMQtEZBGSRAAayrwe5L7dBILI2
qZq7lRKVBfpC1YW+WgZRMTQOqszGNKV2aJwt3RwJWtm6eQsg6PAffzf8XOI34X/0nGnII/KTIuRG
kpjGPb7KsWiiiON+wXn0pH5ssq4uQBO3FiiMTvETikxaoJd09J4B9D5uhg+aJS3duUzjm0/abkj5
GfzO0NCp8AkMKsK6gQhMPHsDNSrYqtonM63kLF3GgPW8Nrl+pjonYojhBpejF4Aq3S+/qY2mR7od
uwObMJYhfXFyJAHvAlchJ0VZg3lOoGWG8kN/giSx6re3gNwv5ostFuETNw25vTIDb09D/2kzapOF
t98SKFVtFGIQVyMGsrlve/c+09EdUur4lCVHZXGFmbRd/rvM2B4KVWczWidrkGpdr39gXa9bG9dY
qaD04xeCZdT25X17x8E9uld/3B+x8oyMeHifQsA01Ye2i5SPwSdY+p4X80DCgEhcajtPS50G9O4v
7nTrF2yveDKtWdXylmczAUwxeiC2l7LtF9ezsc1Q2VtUbuRoKTChqf0pnCNMtNuldmvyfWqJQ+ck
CtJTY+4+vaSQJtEEWfUi5VzacQJb9g8mKJc3tIwvWrdKY5RyOIKj2Uq2ynBNKcEmcIFsp5+HfWRF
5/9MAxjiRLM84VgQwJ5ui/t/ywozAmWRoWMBYYmt00R61J1W62ZWube4bFBYqpbw39JqEg4FXK5J
3C6dzK7Lg/aXajG4WR2MVFX/RsbMHCR9/1ScXNre3nUqdp/Si5189FG2VmNdmNgJ8LvgfUuz+rth
gYaoJ0QYkahcIo4wv2gBZ74U9FB/g2W3/4TIaU5vSdVM9uVl3dtRnZSSF9I5LVR1yL8yAIxjW1Wn
ldxzeK8lxpiHVnUDJFD0NZdiPuuBSFHyXu43NXkcCkE56n954IXv1SYzoFmj3S2WrskF2uDS1Ugt
lgy78iK8UrbyqkgP9UDh3vFNqdMvcy5gM8o4f4xM64nEtkZ0JMOGLyvD2WYNnFcz5SK7bKxWlcMy
ONlqrMDOKLHxcU9FihRR+S08uq9MNRGJ5lIKzPpjQEtb6+Kimb7EYyAsq0s+r35+QU0xClmQqeCs
B3MWb2XwBnngtdPjSey5xYzx8iOm0/D5N0nOC5xgIhAoxRAPqa9ZjbLoK4cNOghlbPN8NbIoq3oq
p1pC4QzbfwVfk7Y01gbEaKUzierOyL4Yd67I+sNTo70Jtm789+Hum743MPyzLoNb6Krx3g1HiMd8
TNCz+Xro2aEvOdRKoEFX093i6Aa14dJN876hBR1ynFbMdOdfQOX2956Dgwxf5axnccxjOJvfh1lX
JPe++V7+ZR/HsgrKpHaWUrm5bK6gQIUxyy6DqbFbeGEg8ifxon+7QplXH09Ij0xcF5h4JS1ubJn8
Novk0Cw2iZe6fJv9C8dCBsJ6pjAbkJuhI0QS3ZmQBSWwUqVPap/6FEDeWbzurz0RZiDT7FmLvx+5
i1tSGh2MbEiB7EmAoBVLgrltyeEvGFNFLaQTH58QOR4RfShNMtFhR7iMhnsDObncTtnnzrlPX3IH
RwvS4kXWOc5bxLbwLWQ+fiz5qhrwI0PrwHxNmRreBWF/TYTJ0xXVxwWbvMHc9iKOJyuFQ0kcvrdt
2uiQmc1v4iQt547AJyctnz3yU+jPCdkzUzMTnQWP9ckOx6cAXBwqyfj0At1gSG9padBIjyPx85WF
If/UgxmWnnIX42k/XimKpAyD5qC7De+ILXgvgsF1xhrGWYJ0nmD99nbVt/+xXKiSMZLZaDo3dt7S
9f0QAqrmj+Ba90PFMx+11LxY3/GdAeKdW2FkkRQ/8uRo3DzHXOXUtO/TkoFomZqEzDCj6oIaF3ZU
UdmDYMy5/ys3MC+42OJbzrwzTHYGSEqcT9R+gcduX1nqDMAGXanp2suYKOhdcr6qIjjr/JuvCOjc
/e7NFNrOYHqXBEXwYX+uV01XPNCegJJ/ol3DnrIrb2vP+y/D4i3QwLxX/796/+e8abPzXhaYCk+o
bGkIbsRWhgJnJGykv2cwUpY2aTN9lg+0c4xy2246wd0hk3teQQr/eJ9G+2ITrFQS15x9YvIxrXgr
GT2wSURCowj0AZQustzn5ml+BQP2tr83USuxJjM+XYnfvr2+xbdm+3gcGIPXpLM5QY4UmynGGkcW
o1PjXVpdo/AaS3dC23XxRr5pLWKOLXuDY0CiB71sbecB4a3S9sPMS7ii/rSkXEOw5anioigtVFJ4
ctuNQGNOYaY1EHv6oKdUZL7Poerw3RIoAjwT8pb5i443vJfrXLn9ZMQkwPgBtBVRai6BKXTEEZod
PFKFaf17q6pWIHdxJhrNToBQE8cRPcsDtqscZuTUxpvS15ij3jzI5C4/84zJQ6Bab5EHbF6FzR9F
8dP/iR5aItTZ4n3HokYC5I3x4/pxIXU2BxzkyM5nxVHdpCXGRuxIJPm6dCL3tTC1xhouGcG8tPIp
mQ2W/jwsZQuc6D9dxzO1WN0EuOav/Wk9+qdyxn7BE+GtVwKrSEwAqnWCMbGnEm/8JK9Tws8pyyXm
fxwkTOu/gPy6l5SEkkbdYpvm3uKeAez0eMCaz/Px7YpdNDrI5++Lx3/W6DYtbq3g5k5v0DLSahvY
hOGgwpTlLehoWHamg9Md7bcDiKTqY2HQN38S5yw8r07Jufv4FnGDEz3B9b7ueB4+sKdPma8rWESi
Y8YIYNCn46RrhE72x62GmoR/uVM8sLN5gc1d9/wlFJ+Q1LoMwRzXpZP1X1Pajd4qqri5B2ZHqhK/
VnXD34+XJTZoo2bsKOhQ3TtKxIzRRMqkuDLTseoxVQzZdd7332rThLFJQtQ/Z/urLtEzCw3d546I
2vd+zoC1n85mGrM2/Vz+1cm5ZlOX2+rQ7Pb5DLjk4HtAHIuWw55qRkSJttdSWvLftQwIEGKSBdSh
jHeXvmbKWLb7PgK2qHTQmVTH7zvacnSzCQ5FKIAPLSSZLM+/7j+7I4ynmrjM+3HBDVX/fSStaBAW
vvZHBa9a3UXbHB8jBBVeQWdP4F1fS0j1m6OQyRnWU+Ru30pYLVnBt0utuFPiOw1Wl1oHk9uOcUNR
0/VpyStxwA1xAx95IVKDPqiyCASh4EFcDgWa7gWZhj1jh4Wj5bAsD30obJhzAC+HkSnpjfCN6WjR
rVy3zfTY/eboFwj7//EnTrh/qfMd2sHsamS27uBkDS6yfCpttQcCAg8URUQcS8E+Lrjgba0inc4T
FZ00rWl4vMu9A7mpv13Ai8U+Wv18yWPgKAdtg389VbTYJCSWmsO7OE5WIFoGUwRp7TgRN1nCykVN
Mk0utIMXGHnDOtsMpQWa73lDVBzEYhpjWdTm64O5eata94P3zWGSm897vL4xBkJIwf5QIrdpVo7U
0YMlWI0gn8Sr9+eFpUgj+8UjvQzIFYwjs/wsEd7vDSLkS6I0BJotl144xv3q9LfOy3pONXeEMgVA
Mo0syxhH1EzrQ1FkDeePAQ2JwqjJDJW/8LNDW++GhueGYL2ylhdpWACE3fprEEUiR8iZKYauuEY3
b04FlGuOz499b1KGsvDMNkJTOfOifAhJBusE7ao2n0w4NQYnvvsPgTGkmp1pMMgZk2Hnz46EYv35
QLDU7pp5vwYJLCB9SZHNR1r4tKItPdgcuCcX0zeLWk+tPUVSHWVqGpqq1NvJn7Ze/bbcywDJRwZG
1uH6W/0ocIF9IlutgXyFkm/tknQ0NJC7U/p6hcj6+ng8KF9Ttux9rYXHFQL34MqvrM/YOU3bt/cx
HOfymqbUur9O7s3Sep9AFnp1ZxgJV9hqsA2r5rk+ADJeGojdEqpSrSgNRNci3B0fbyRXjnu4N9d4
2/6xihh75aMqSblTfTsiy2W0zr3uLDrLWILdbg9MhxounStROpdkmdZQ2H3Mu063GvaXuynqZRhl
RmeNZXgWQ7TznrKXU8oa8RTlS2p1mI9PHD4QWiKI1JzCS7OTsZXr2BMrakkhl7Apv2il6qKaIVP7
cTuWkOQlwRRGhQcG0m969EEbajyurHHrJr+0bkrClw3DgStHxYeTwoRK9uH/gSQ2KW+av9zIrQ9d
qGI6aJ+a2S6BYcgOUAUjKZOaImWvvkYsbaz0JzYHy62yHSClqlylumUe8bAkoeekPVNws2C4IHsN
gUhxc9zurftaYVivH3df1pRdHotUHFBMOyreWDPa1C1ORxLHVyJKh6GPjaan0O4YKtdCRW5tDAW6
I88SQ8xdLzdbfJ5wlp72AyoZChN2N0e0qT9HWaqZsOnptmhKWzKAm9IQ+KR9tPuKqJgmzojvUiIw
0WTItkBPuV3pEUW2XBY4wRP/lseWmgG/6Xq9SY4T3x2rLN2jMLHnwhh93nZMooCgL3WySGYVsOL6
dW2CMccMmUshuIp3pzyyCzEqxldGpCj5p3knGNfN9Kn2ozBwad7ARG8sP5JR6M9CmbMQTjQgDyGK
FUwFvoPeCfG8bXdoW0PyhabZnlUgo8Hj8dskujkXqcni0T8p29U0Qc6H29HVfEPIWmmy6H5/lAFD
jNkRmNOANDz2ZQrDS3nC/E4is1GF3Xj2o0jU4L5Lj7WBaKS8+4fKbAHIiyitNGqZEhHbzzIeYuiU
+WI+vYOtG4o7q3RqR+BLR8KMZa7wL8dOTWzd4E4YSeSITUIGbpiMBO35wHTS6iBgExN6xOzVmYvN
hV848CrGE3k8oVEKl8ki2jngaDbhY6kEqNSJl5xcuw5WU0jPQa1hHItUJBG5ydcWsbmriVLcxIFo
VqNTnXF4pXYeNFwl6mo98syXNjg29Tu3wCjv8JzvECQjUKyPOVXXRvrXlDrhZ3uF4ndQz4SDHK0L
KgXnjuIVr2zwMPeKomVckWj6pFfUwFHbY4qNopEb3ASbD/Imwi4jkYA0zhjGHfulKF6sVZiukTpq
H1ARAYJaHuRvTXg3ULGxb9AQxAdvv3Uk15HSxWCfjjPiXOQ1R1imaRh5NbtrTjWWHWGfAGhAZnlq
fIhl7qQ+THcG6wUNNQN/8oSnWCGyJ5+rmdFd2eHxctvLfwyhv5JnqyrO8xOFLeZLcIW3qu6v37sp
ECvByfd2JkjsGz6aTbMhn8L3OlwfwkfL1Eqnq/Xu3Tdmt7zzEH+Qua/X2Nh8D9JlTjNQdT5hlFkn
cc57WzKGjrBapbajmYCrAIZUMEyKMFZi2nn5FPgyQj2VIU7teOo8n4LH6uKC47gQ+k6Sp7/WCJK2
Yr2pI5KXwYh6gWIjO2scgl+9Ma9COq3plUE1B22zqQNoambtjliCXylEkMGOUkS9TGJW8DjKV+VJ
k2+KJiXAbd89tIQC7Hl5G9ZJQ2MgBqrCzJDaSHVvMpoXa8rOEuJLDezWbKKSVOeZmjsGsFIVRBM6
7XZSy87y5C5F7+WHj3YqnXtUNEsQacg6wSWC2SiPYbX+S0/d4Zc839zx5ySqQPSd6qcjpAcKNezW
XyTCHZIaJco5V3K3Yd/Fx4PD4Z4Wg84VL5pDjdivztTS1xSRUmNuILjo8cykomvguFkyfz9tv5xo
/pa1c0HSJ3vZa02XXSs7Z2RYnDe00jzR0oW11jvL9kzcW6KIHQKt0BYZyMH58syt80e+tk/56YYO
seZls4yRCQxEjwwd5GGMmU/SNRkpR3Byoef+ARKvRreRcwg5g619bikB1z9h5ZvdrHd3aoKTv59F
OfuBrqMAqL67jwgW+1nFrVTw6md955twKV6s6K7trqMO7D2AsICAa3BnEZUuQeW2JLAmiZp0VjX8
cyAqZXuVCvzyUIbHB5/z5406Xw4AQXwWbHsfhq8J3EI6d8pAUesYJaXDdmDUfK6Sk1YEsAmkwdF4
iF0Aa4vKRNW77zcMNU9uiCWP2RoO7RqjFmNGvh01W99lbdnTPpDAUddM+PjDJHrbrgarALEU90+M
M/TaRjgqNHumc5CrRObq+pwBSLK4F23pzweumZBqD7bQVKRe61WlWQ1JOH88Oub8cRvn5r+BU6y7
SY5pw77pQoYh7Br1GbwcUC/8/6YX+MSoSdtM8t8r4+77a/jsgEkJTK9D4A74oqg28bL9YK7l1ar5
whHMm6Kb0QDbhNtjDiOwL1/i4/eA1JSOI8+WycF+1Tu9GN7zwXuG19ORB5xO3N/eGlPxP+kwUdss
4xE88A+NRwwUEp6DYEBXYzrcn/QPbl2u+gjlno+CYdycXBIxpBbvZcoeqc1ipaZYDrnAWnpp2Vf5
5OVZVYEVQJLmCSW9zkxklIxQZkWta/Dq4A23MaDPxOti3EXyQQi9MCzGB3W1FuvO5QPHUMth7Lcc
SBJVAbC2jAf429XPFgkHdJL9QAjkfJR2QuJBMM7Wr0LnYe74yUcg1VpT8LFV5TQNU4jOeCAbRfSw
kiQJJcMFred6gfnicJV+NU3Bc2BGGwonzk/I58iCdY4ASET8gyiJ7ApkVW48MIsU+3fthjKau+/J
RbUY/UZA1OIlgUV6rVaOtcyQHishL3umzGgRrkGpgzbTO4oqnNMbw5hR8q4tdcr6V+s4jzInt6Lr
fJeWf/2n4QQYPYX7XDNpg9aqOZSCy06hRkW5EMAIwmuabsYe2DmZAr58qLAzYIkL5bt752/vzAVL
/EoMBBCknNpYAXoPhdQUUMlvLfXH07YQO6mRFPbIYC/oKeuH61owV9UA308sdtfNRoNCIc+jIjIn
zX0ECo4IvaCyvPni9BOYNipGwp0jYHimo5WeH/+F1Rf51neJ8HM113FbxTgRNB+OGv1KOugdbG79
NZLx+GxmKDFvVNU+SY+yxpTf8E4T1Y1ZeQiGpFTWH3Et30xXGK6Iy10lrEaNb5bPuFeF70Q/5c3H
jNDRR8gi2AAx2xJLvhACTW364n5MJW0Vt4/ek6z2vPijNCUWB41eRSG44uYcSXYxwX4eME5+zBYO
NsYYs3HMktdm/U++RtyACzlV957z+J1VHVV9/+ggBCAGgQHsAr5xs/gddu3ab3D5fbVGN0Cnp/H6
P+YRRxSIuVvyp9YQl5yg//2dGpKspA8PDbMeZGSVFL66N8mdyBI4TIVj94K92VMpg9pDwB6Epni9
VDHjqq39zw2PausUoKuT82QKUqlr9su8VIIvWUWTL9tTRJnY2LfzfL6oBCe89CDdHX69591gZGIq
4GAk7gIYgjg+ZYRXZy7P260zOlQF/hV8FW0G5Oqr/L93FMB9SPXUC6jj/iUFs0OPAxCXmhMFLqcD
ddckH6j1h6800qmOqMqjFX1v56ICyi3bAqKbp8FA8D2WN3qCC4EO4JSP2oqFEPC+FxMkZCVuZgYB
DqUfilpHM0PCXDj6+0ig6SuaaQtc4E8q5g0nRvS5a01E0gtv641lSz4zibzgSjgxyW/pDE4i5FjU
huC+gORpAL2HPT+WrbfK+AdjcMA7dH8I33HYH3vptX39lTkjNSiSaO5xJq3VnyDg7hNq2Yx1Zi+r
EXHHDd01+37gFpcesQmpO3Z2xsBHEc/SY1tLYschGd9r+3EUIZsMBz8PP9EZmimDTP51cXv5Shz2
NKa2xIUMOrk0JW3BBSPWJasXbTDj7NQcyii6dtPkKX9jiQV9a20MjewGGeuq63xXiV6zFZuJpKRv
Jw1HQVTWd//KbtDSyYZvKOqtce3fAg3Pff2budS/hxyFuCVHVdTTqL9NP8rl4/rXfVcjfn76pB6Z
yHt6vpYUYa82DPRDJPbkky8bok0xstr1LvE+ypRY2fLVbHDoo1qq5UgsqYgJR6WW+6SshD0vPmzr
GNOmUd/UY5uJG3acjMNQthxwnQwfie3ia7V+fHMQhQniQwdJ5rfmTBTSZ6y7Qg7SZ2rFIlZcae6t
Pq38A9U812FT1OhZjAXiE/MUO0VGa2gKWGGLrqeTBF80BgPKXk//hY2hTaBlmYacNL1Va5qy7Aqa
X6lBWPxySOPIv37loRybl1I3YrxO6SuiH0m09KI/6/m3CX1rKh9wpTzy6wCkJuI1WZOT4UOJnrkM
1ztummo/jNcWl38nS0Kz0puzHNKGkji1R5BaZN48hMNrimPXinnG+ifHS3BuRrUUMq+EanZhWUAP
NSv8nqxs8Kw1HooMoTGUVBcpzFh8X1xYE3SZDk6uuMnt1e25J5oS/NKBI3gwwA0T+BsMROHMNq6h
Prv0kji1k8DvdZiGj4Bf+RBjHlUyOHUB9I7ZOg+tXdujRElLRFN+xS6FLDWX+m0qydF+O6k5iCTE
nCUJ7kQLiiZNh0AzkMvcsuNvBCCD/kqW/9OAA25v7+/zv/lJ1HbsChzJb0mMMabiRpQddSsnWKzT
UT57lkXp1CnJ9jjr6iX4nM3S2Z1CIGvNt9DOHUGDRgk6wI6vE5Bhmq/lk4bDnro27RSkkMWFUFKK
dFhDfULpVRKUU1BgU+ly/Rz9gO0hDMIXAR/HLUhPWBa8R6Ziej30byu/ILRlW7WoZ9gtSF6IWzso
D59/e0xpJvSn2wF+tJbYy7624Mt+3e7BOsfqujORlfvRUWJ33g1UHRE79a8wDoMxA9cgOBTtN+iL
Lmq5yaATrlHKSt2CWt6UvDOu5OVnVPhR0ptfghUNrezV09PiL0U2IbRU/71pMcR6TK4rABQtQqup
FVbRqEw4XKh51mz6T12n7TipYMmksfCiU53Fm6rv9jh4PIZuGXI9SUHWC1/MfxKqVaKD5ccxxpQ7
N+drjsPXSc9Idibo67q4QihuOvt8uok+t8bAzV0xL4RDC1vZ4FjmaqIcIsXpZBYI52sJCIsT9BAE
foLkfuMm36KbK8+/aowiC6E0cOmLtiIGJ0DISc7C0stZZUut63IA7naxZZ87NW1P57bjJtiWv3dc
2X6/x6qNV8m6BvmCSlIkZxXT1nRHCphO4u/hSzCsK8xeFySZPsJYoNlknV9gmzdUk/CMLKXEU4BV
1fHF1bskNlDehDqO6gY4Jk6PqXdKYghScJk8XZYIauDmX/INLYiifoTSbCVK6qHCGi9371/y2b3I
TPvLMpTuVTVRJs7o9FDvu9dh122ydaoCVG2ZDMrN4D3P+orWG/JN9TFQ2rrly6F+ZZd+HV20laHu
XlfSDpB1f/GhSUX5XvlmCazclYTqmas/hOqNHCem7jC5Y2QvwzWK3QHPW5gOFiYQzUT4JkWrfGoo
V0buxlXYeUWNTfE6P3bf2UzjlIeiulnZHP61DvWrMyCSxzBnLK/KDrXVvRifY3AZZBtruwvAaCJm
+AUv2caFZ61PPwYjrKa3TGUgMgJ9PPb5kk7pQVLRGiCCfsmRt3bk5kx1+rYsxeMZwoX/9CjmbsVW
ML1t5NOWW59R81lGUOlofCC/J/+Nwq9+JbNwwYepscx/hlQ4mEGAzoW5gT/ML/lHbbbctr8Qr+QL
B6Ma/tCcwfV3xUnJPicrw+u2i6K51SjYrfUJYYs3QG5iZ6/yxbQlfwkWFAjfgGUWSdW09TKgFhfa
lT7zGdjHLtGGk5ERf7hrBCGjfdF73vXKQSTJncdznLF9UCUKZ9brPh5ftzRlCFaTyePhwI6/+Gqk
ImvVATA7Czx3lKpMxZJwyow9dQDpAGMw22SEhdjEw4vRvq2XLmeYQmUv7jynX54eZrJxjSGRiYw/
d4ctwqxh5V65PbLt/AxnZo+0D1PTwi/kAStkvLDqYiAGr3rS/jRd+FfTN1yGB37VhsaH9iLdOWAQ
V8jQXNHDBW8UlYvHSC1WGAqkc058OxeNq2EvUlggsowuBBDS5QwCXz7moWuMEeCfPJSM/K0s6eUQ
6j9TyZVC5Qk9phe7t7rehu3UW4W+S9BgWLYE0d0Car27PH2AWU0ygqSGR87iCXc8URVRUkfEnVky
E9HWddx1Plf9IjViOH97cETAcWOZLJJ2GWYCDBujkEn4AKhnOvhF03qwaG7fYdd8DYjk62wcWXcH
BRoYxTc8Rl5A2hfHbYSBnZkWMQRs4LQB4Mc5ENWArvN66FPfVwmUoe/a6ur7pvN2ew+QbaRG8Yqw
tFXBydwUJkRUY7YGwxabFERKJz3prkRt76mJs2dgWY4Smx+YD7ZmknDGLE1/8/1lHDpKNyzl6nDY
4cWNwCDb1zitkZr4CYxKVZ0qGgNdojjsY6GII3sRBOh1q1BhwAh1lPaI30zpO1tAYYawgMu7mkdC
PnXVdLHgek/rggIDXeN6TqpYvuZ0TxY+GI5AGhkhNtKbpWs2a+XoT5X/etXfQIWVO+p/lgqDPd2Y
yWmE7TNsHgIRVfKEc1Qxc649xSatAIl+0huGEorisHv3JkUQYRYqvUeVxFAtmIgjiVpw4mUQWMPu
7TKhJs1Yka9m6wAEUVVk2FV5/3VFZ3/IEZ5EAYHKhvGZEi14X7SQmFbo9QoKRqqmHGLVKrJw0CJz
n97tsqJjFELfgjxi/R2Px5JE2xr18VojH4InE326bV0ahdLbtE+inynpimacGcm1ArLxQS+n6kMJ
7HAVYO3WrbAFSdYN1AGMLF4E9ShXmhnH+99ARfauaS5FWonhReDMN52WxNxilCnuk/J0kyXc3hsu
aBE/qAxRihykUa6BnGMHVhMInYkovMO8D6IIhF9KqGo0qIuKY+dyhMcCQusNIyXZu92VQnF8H0y7
OCtpyC9uxFFqYq+Z2u+01HWxsEdCkgT4qiJCjKr5GXjKnpApQktfv3CSbuorbXcYl9ArQV4hROX+
8qJUXSJYayCJZDIMSQp7908eIaD/xHA4IbpFXXSKkM9sQUVaoYV/xRC5bvMQh7qg8kEmdWCTfJUK
q2NC/tRLnq76AzNa4ibJtXxla/U4gw7BcKCZ5Gxi+kFa1tKaIJsCNa1nTlVFKiXeEE9+ZXfXOYe8
F72cwoK+csZpozLh1nrl5og5dcdqTcLNUOtlSnyRH15X58Z4zJ6l/klegFkyWeluxEnndEZGGpQG
HiXd/RtLea2aST2pmS0R0w5eZFCKjFlotOtzPKjSabKbqFBFl5I6trIvuhc/zXEAPrOCOPWNYGI2
HwM0OJJuU7cnHo0znKax706jogzMskD8s/45tO7I77TIBxwLf6sci3V/WsKP2ampDQamJLaoFaf6
z3AQeAUeLUPZIcxfqX2pCKPLWpJr3izERClHJIeMFpkO2ECakCxkCr/NsutGGY8m+1DVJvd5LG4w
HLRB0BsQ14FIhfZ9Q3YHZ/+FYy6+Lq19xqYjpJw1GgouiTFUqhDDuqY3zvDaxwsdl9Xn5Amp6WIi
JCDNZzS6pf3loyOZKLmslq1XQGLkarakfEIMQkyFzowi3YqTrh90ERHeAEWhiDpBci+61l+kXG/B
HTRN4mMNiKnoeVzroapWGU93KWfrHete3tZEMacoIjNcbX0GnXrNL1hs6Cd8gkhqpkQFsaedD2rb
L0p3GcNZItkUdi87nm4AAM0G1kJ1yrqEvXkh4++TlT8rjzn1jv31nqMWXjJspvt+TbsePtmPOzeO
bQsH1e+dzNMdmbkHkuT02MoUh9Qxt16wEox/EimW9foIJzV/5+3aFz8JSW6teJ4XyGagLebUs1Lh
PPUIYI5uQUvfpJ1Z0tBJlaxXhnZE5BzfdWSA/ZSoDI4Jg30lC0qM+RVku05/qgGnpi2q+0TNNa/j
1ytPEi1gRip4JLoADkhsVbvretphGmczgxOMi2NsOo7IwSaKhySe2fgw4g92IXJk9ZUso2TiH7z/
tUl6uaTfhF4aCb7IDxMJ+nu6vGRZO6Qq1YgMuaTc3b0e+a7RW2iGplgMP9iLm+jNvlLZM0KNoQYD
vOH2UrVCnaG7Op1ZsPvPT19yVSntVuDEOKesy1arWKyeBoRCBvbPrzYGhKtFrbLPpE5pYY3sZjFq
fYxvRg6aZ8JsJAQ/liQ7OBRZTMW2xhkXMW4YNEp7gMw7WTHJ8jk4eK4Ct5+y6+jKMzLI3Nw8i/PE
u/FSC2ToRQVNG/cNqXNIZILUFDZfFLMLV56IKsOXVZECi6WPsvfGsuw4EUf4KKwPfGARvDgiiA1t
UyLWrpMApE97uY/Q2lK4VH0XYi3WVV7gHpcl8ZgXnZBlIeETTxKm/AsmXrMtMuXW20TvBZuUuD1D
rrWoWHzfiuqxRid6IeWga1Al0oUG6xN5TS/rOBPcOuPRSHe/m/1aKQOPlme2X6mz3RZ+wtUzpX0O
69ZofTdBgHjmMmO7PAjhhLgZpRMMBMDktTVm/yCFPvc8AUzy51g5e9i8gqHxjUOoJPrz4DwIrR65
2teDAWilA0zKEcCXp7RT1yoFSBTQOSKf0Q/QFNmQXt/ADp7zzl1P+pDuivu5e7fpznVrhCryoSaz
r+3vYR3v6dIg37GMQFuEtX/mn1uL0aIuvJzhDZ9PSm1Mx4+3YVczRx9Th/UfEXmsN3v7wE6gps67
aafBvv3gczyedz4SF98xsqyYXhg3ByOAkuBUQ/PQQ2E34m48yDmDnQpMT/cINjW3hj3gm93K4+Hi
cA9uodVaH8Kq4+Oilxm/yH/QzITLQMbrL6I3HVnyKM9wDElbKxxQ5yhvWLlRG0SE7oLwk3tVf/0x
EOqA69TSZksfnSDnyXGHtnGQLzJ6D1gPKRHdSORwGs7+gtSvsY4XFm851H2GXAivoWqf0thsUgse
cCe3MRSqJp7Hwb3nhScQODoA4mCpS8kxulgsrnhZ/S+vFgThbycxdSGlgp8cwEUimNaM+x46rbrL
A6NdBochG56qV0HRAMn5ziP/DpFG5JFzkpIsZAqmtvSKRuKawsd4mBkc3CMeVRnX+05VmKgj9JGL
Bdy/tvN0K3TJTH4qisfq38LJYpbNhCF8lBbma8zQ89gLdnL2t9fj2M6uNiuuXhrMzT7s+Dj3sqHh
Hu8q8XF4xucwf0NBFr9ZUkqyWSuPqZtRknBESB1tFn0I3DM8Mxq5h5FAohd8N658KkqbCEC7VCin
jtuYfC43E9WXJ0V3Xe1AGyn689Uo1F2cqMr1V1DJocIkPY/GOMItYStrF+8+4dvU2kXhyHbJ75fS
tGIfXIl+NYXg2lWuJMO5qXgx5wmio5m7/XAB8RGE6DAIFC6BJtW63tsKyRy3zleNXTNBAQB9bqY2
rOR6UZipiqB3RmI0GIXrwN1Ikm3b9FPC4pXucsTRZcM7WV5xk+9h9qnhanZIc1nLPqNS1bhL3qkT
agFysNnpa8FXQ/jX52uJpX0CXyzKG4j7J/xMEsEHf/PnsXw3NEfnWcF8uIzi0drKF1YLzuKxBiFn
D8ylQAS9QsdyJBreUk7jEQHgPjNkLsuuQQhdOoZtxMvICP1WVKpefw8mR7n+6TOCjGR48TOnwSoh
oBMfWUHXsnfZZtvZWSQ2mOK5P2aK8Ib6cyck4LmAft0GUIHoN+pp/IRlJI8z1BojMyo44Cxq9rhf
0w8PsDtDJmxovT3Nho+mZCO+halYuzRYlGlDvs5yuAPbXF+Zx/KvhyufzK4Nx44G9Qx/MeGPNYCf
cUpzNQ1KU47cGSEZUTdEUWi3mipcy+szi/y2fm4kgVpYrL2G3oIYKNJ/s8yK5oPNPgEDDd6vW1r3
oBQ33mui1QKgy+z2E43UGpxgrDlP39KM20i3nNlvIpkzmcc/Rv4dqqOADopurPmpI68Y4mYxyjzy
YCXBw3YM6IGr7CriB7lM5PWFm/Vshm+GrFBSbS75P8J5Zo1oYKOl8YrxOOFDXgWWgREvDYPyf4wS
N8isZzGFUAc7Hn6MoNTellnVh+jPSP49+j5CBI3TvOQRL1xIxKW1On3SlCVXOB7Afj70ps0pF7FV
BwQJG4kyhNi8hv0lDMGVtM7Qkw6NsP5lWDnmsruGdAylw+4oi2aherAgcV6OroDbyljZKGH+uhrd
WEcdPW2GTGlyeFLJzWI7JN6Bf19zPN+y/FSHS3BgZypT9q1ciPGFkC7r++LM3BlFoHnxx1CZVRn+
T+pGxL1whTXUUMxaZyQ/CmV2jVnVh+lcSjoZU8qwoLz97iZJbMePlzM/4ZkPmlXT3JXej+UDZKL/
oHddnObngno3HC9obzbncOY2apeK16uwIKSDVs57TefTEECDSzwZyZUnpnI+P4UC0LpY+3cWEQNZ
lvu62RB9SmGSqnb2Om2iAles9QHQcwbHnGunhgHyoffw4TGM5Y0WvoCosrNyHn2S0aiXZglo/ryp
u+M2AuIsf8ey7CENSbgsb3N7p0yS3MfAe8O3H4558Z3aRHejMhbfvbcwpB0KnYVW/YLchhgVu07S
4elRjcdBdoxwT78h8bJ/jqUsV1nLBUyoWR6UG9bR1Y4PD3vMBZJeWWAWEPqKhB4RXE9MZFPKPNLr
WAasCKVghHV6+r7qzhiH/56z8z70wi0GSzBKEQeBH3Lseap8yVwVWCeVfTF0pRnKyU/e0j5uLllv
YXKbHvynT+o7rYNcxtsEn/u1xv9vkE+0zsqrNY8D38FthE2ZIoFrT5XmdNzn0ODNSipJPsfiW7qq
pCcLafY6HYvYX/fVz6avSNVDDqz75A4dt+iikDtEXY3SD7TB9u/BGVJNGgkYzI8aS2n580ioyg6O
s6o0Caog1BI0VTxbGD3vI95ScqFaGMpudvzUXXqskUvVL/33NJMSgvo+KVIj6O3xA7yllxWdgV90
u2e1Tsk2FGQu7X3kyt0GqXZiR/29XQsuXh3LmsgZ6nRnaSNqzcR9TxgIj58is51YV4Ltg5/D3Tb+
x0smjz3yBNkZVwKamAFAG2nrWpUnbMvuC6NoNXMl7kndoP429WY1XI65D75I0ktTzYMKQqB5pP2o
nwcogX92s/iIhD/CIcekYfFFJ8tKStKl8Rg8Ju90vf5mVOSWVKvtZxJF2L4Ze6DAU20/8PmjDzpU
9FQRawL36ktlM/yp/QzfCBECamfunl6gQ9oSUqV+/I6pB86lT1SPM2xg0ZwpsF1P5W+xFBHdvQLi
8zHZApOZfG9ZJS6SzICDP+CnmmMzUFgOTsM1dbezUfiPEL+np35ChFAN8AojamVIPHBxV9aw4u2/
qys4hbwvU4TNS5LJlvZprfM3z5peepzLD8mqgGfOJbJstgU0e+MRKf0M21iv+OhU8vajnymulUC6
xVOoGb6IHJ+MCMs8FmkInsNRApcoCb2F0htEPHGaQfIxIiwlfemawIAKQsiO7s1ZRPYsWMqZl9qO
XAgwXs6Hpzs7QJVVW75PhPD/S8nF1Zg7evvACyfnoa3vFp8LeL0A3/4vKn5gRsw5yHRWehzEheQt
pvkY0u9xX25+EujS0JRr+3j1j0Ry9hdZ6yCgQ0Y0s/JhmM+W2ICaqyzus11ab2DP6EL8G/anc6xx
SeWhe8ph4CNeNT1pGBu+BsMjRjTeBfklgfEIBhYpitSUDtI1waxusAmcQfROFC71DyZ1THmyzoS0
rAcrmP0MdfkGw8N0Ydgdqm+QHtCH/XzJJ/y54+/M0WWlE8ii7ZhamU5A0yhd8c9Mwlmipn2XZRzM
ZVW+4JzYyp4mHFk1nZIJAG90nAvp32lf7FlXlDSJ++RKoz2NIbE4jImyT/XX3u2gmZKRRWIt5G11
miZLY+oRfXfdadcJ8yVIoLbKBPXCN6C4IvKs/6z7/lYfrCC91qJuFZdheGTDP/ygDsUVsi9cpPT/
dJUssTsy88EClf75yLc9xT3ziyBvsnX7Zhqy/B+thF2+1lZIr5Ji5eU5NjM3s7dpZ7UPNh+O+Woz
GhSfuSojuHwP3zTDmKPKdLCuLXPqtu4tds4+uCUscVX22pA4Ofa/BLcRNlgAfSi+QpE6pk2PMIib
uxKZSePaUt0X1wZkt6phJ863+dX6HwMxypiIaR8YkdbVLWpiyHr1vBNA/tunk7qEZaZLGOAG7gWs
/TFmAEAWUMay44f8IKj7Iheju0Ms2+u+8/3Uj02rC6WU2YJIFdCa2OxxhYNRll5mqkE5QhiPRNuo
sytBloyHdKDE+GumMYT1h7+IKLRYSlprJlgd8zizGudCB0sRhsX9QLU0l53Yb9J6xTwwnU1na2wZ
hPLtVEexKzzSLM6SBBo5ku2PsNnDdtdHESGAYg+IytvLKcWooKQJj5GXMEL6baGDoi1nCIBfH5Vt
XPDf+2IU7s8kTPN24ZxCTuP9zalhVgxy0BbCZxYhIeK87+oB31kV3H1wsZc7RO5avNIIaJ4fpBPJ
66Wv9kqe76Y/t8lJ0RfO/OnGbCzL9b4xVSR41sbcOxXzbN5nE/03SxgcLeovyX5syJNd8cmrboQU
6XvdkU23lgYvu2zL3oIZsg6jPYzRwDAa3Fp+sB3ESqqv5jKlr9ZjqkutGy1eG7k5XSN95pXU89Yg
jjJQ6a28QuHEU0HvZBJe8tOW70ABdOGfPdccxqx3/eS+qtJ4E3jxVYIxnJGu4erxJXs+80ccCXvN
3yNXvHswuKPFa3tfbILoo8IoN41YYBY0vX+AZ9Ig6h6uxv8/GDJY5UZUYZ+9Iq7XmtGpS8mqP9i7
UhI0KehiJUi6UMXwu0md23+h0WsP43Rfsh+pfoUa6vUxVcPjO5umejf84DtMsJF+bx02iqGFCtp1
CMAkXsJ3yXj3An+INzJegmAH8me2/oasNi6skGvhcgJe1HW3rz77aGKqhYkLTCcMtCbsUtgeFe4w
nmo+g6owB2wcmdNb7KF2kRoOXEbBqWzTXRzbOjIZOFNoHm0sp+v9vjEPbODRotZygrWGZ13fTRff
2bwfT10IKhusdHccHD8NSGCeT6WcaTjCfnpcnSOiWZvDBuNZRwf0PRtoNf3TyXu7nwakqUjVzUVC
rs8sUSAtOe4VwrMpjRCSn8U5IopMbNKne2Il54ih7Xo4wB1kub/eSt/6l6z3xaOasxmSeQ8jGuJK
lw67tV1HZVHmmKFfj1ej0O5URKDYQwoTa86jFyT8fZ1CPuDD1Pk8QQ3OPZJbb70gH/imQjTI+fxx
/F7JBYbjp3hlXX953LrG2QccA+P2uA622d3+Isxgp7lyVqhmtoE0TjgxEAJToABxLWJP5iJiDQiv
WxxZe7f5U7MmL3tFzf0hL6fHrlEDu1VoJnJE/P5lz9c9/1AGmGcDa+GNCdxM66W3PhUXydTa2Xd2
8tFAWDTcsMv8hSayTDl5pnwXIigKs6L2fqT/HS/cK9EhUrztHLjdhLjgB7bC5EbNskt4yU7jRv1b
QW82dLafWApNfCLL8Zmqvwg9TwbmcNEN0EkvtdmjJTxjzJBIxTu/qjLnANwbJubxc31w8I4hFFtU
vn3ZOmhyC3mi+2kEDfa3HaG7C2QFw6e/lC60SvGODSh9IX9ZHi+x0Kt5HG4S6Hf0cFlq28hXtpk1
hFlzUBN05bMdgJb+ZOrHyeT7k5UvChAhxbTqptUr/2X9SUnPlMMJcJgLlLr5BQlywqHW2Vmj5Hmq
jwQR0vVB2cyt+kEQ4aoj5f2DZJStODVcu9mhJx53zCkld5CSWCOcuNcIsLjf8Vw3D2Fr9/L66jA+
sGXZ33yc5Z826ixwipqDzvPcErQlOqBziQL9mx1PDiTFQjtghvOpzeH22mZjOf7k4sXd4/ZXJAxE
q/2MqY+s9kjM6wifSWWNTyFy5GQhhTzVbNo1VpQGtlaxK2DaZq15/B7ThObPsliUmYrCEv0pWEj8
+Q0T+72PPc3DgQWjNRwwl7DxpW5CnrvohJhkBIzzYVlNvknhjSYF1RFU/iliJ1CXQs9v2Gy+ovnY
ZmnylS3ww0jG2pOX4GI2D4HJiHfq4orT2oyrzwCU5TmVAwOXoS0XGk0j/uSF9j9BLVKGOOOHmuVj
kICj8JECG3RqXP7rZzmSg4nykcs6uin5UhuveW/Lhiv436Uu/26TBm2Keo44ZWY4V72oYUFJ9xtk
7KNkBPIyGg0FSBleA7gmze6wfzraXkvuKq3ssgJUG6AE5l3mwZTc4733DQzpVx7Sn3ZELdF7+wWA
lnyD/FlsIR0E9jLnm7zTrywhT/TQ65/pYc+7kbBSHFJZeEQAolXNvLjMZsQ6LZBWK4ipMjBRGLw6
OzLdHq0V992E1yFrloglTiC2ghOUHczkYLc/iifUeRnmixW8CCU7syfzA+0uM14afaw13AZjNnaC
3NyKfvUHhXBC+2lFQsOWBh3Rhx6nFfw91VIKj0aRU+rLuhSXY9znBwd/iIBoiplyeM1QiTu8yZ0u
5wAYnST8XKbOZEhLxFNTA8/jZ2HATM5849CMMdU/Vgg+C4wiYiyq7UQRCwFDzDJhEvqDwxInhNka
n5Q3i9l3fbZdGXe/InZu762G+KYKwimTu/WdSPQyvM2HZ5/IJD6JAjgKS0LVmOFeYYVGHawS358x
aTt6v7QagmfZdrfMYz6dSZYFuJSXJ7cph8RggMfTPW7yYZ0EthvSd8KDz6cdZIu7/1IC0/f0aGmS
WiIojL8eA6KxVfd4Ps2cbon7+1MKEaE3GRbvpigoruFhh7gn9rG3YgsA3VI2dZlT5yUFVqB3lCUL
3CaXDCw8eVelOFDUdJv8TKdhd+9qeKRYWUNLfOI7mmgVnHXdoLK/p72iY0CjR+i+7ZsiAruqhl7W
hdHwkSAfw8Q1pQF9o+jNh1g4m7pL/a2PID1mlO3OwBlcwW3gljbjNS5lqW1cTriM6w2iVNDD/i3V
sipSWbgEVT9D8LJluwxjoe9PGpNK9OwdI/0ws5la8voVQguSNLFiTl8nzJ/3tKOOHyX7DLn08MMW
SyB/+eFHwRDHY6+/pKplt224VU2qwwoUaovEcjccEFAUI+ab8Uvh7vtdFPsREoxQBO5JZPM6iUbv
rXNiHDWptCXkVlELzOgu2cwJQJs3/s902SoqytlVP5PwLWSDFhLMgUnf8rGETx7U4kCqaOunFS5A
81ovhjiWR/4M1Pgz2BXLYheYVq7MlVZQ43rDM1PoNw5V2wEGhghVg+rS4TOqIflDl/aEpZ9CIiJX
V/cdTVkemI7oRu5diqmx1ZWWfiIdP+rhEzO8izsMDXYhhCDdXImudxvvzk3Rj5tiPa5FWIcYN+3e
EuY9/5BsrkUz7bjt6FcJMkiX+GZVpFQ5EqgbhT/xL5czLx+fhkbUpwK0LhFuceZOwRQLKjR26U0+
1JBM4VuDGbxFnn99WysM3l8fDnnnqBsLRGUGKdJBbbBWwrJv3n4+qnpJUNVwYKYqwbCbmzj7ZJHk
rCbBxTXveUms1iuVnMBWeuCAqWUwHu1JFu9e2TZDd0z5yrRdX2c6+SlrEX8NZwkDtKnGaSKc3cLe
gRe47MsMj8hSgwI8EJE6iYEyzhMqw3s8jfLMO6Jj3fAVlPfJSyzNkLkiQ61j7M8nAaL9og0NAb2J
CDkcfYwiXhvfvqPeQqWjkgdBxlR/SNAySt4Vkh3F8U/Y/lnTwU/sQ1v7tJhFB5TmZlxG16+BGfk5
lXkADz43gCnUfxiCa+dGp4rAVjr0xdonoOUOYsCJdGSPGPfxEH2Fa+EWILGaSEgMLOFMA3+ozxXC
gKnCe+ui7BvwW27VCr8TqrMELZjMtra3P07LUbML94lVFZP+zbAFd/i1QQ4tDNYghxfoDzwHYWar
QxGhe99c8w+vaF+OTLpog5L0f3tMlOKVgKmYdE6seMO5dP6+CEr3PCWIx90jRGgdnTK0dojg4gKx
2qU3QxLFVF5RmrqJttsUckNe3xfYeCtve4S8Fb22zxYsmP3A/FV2XWyiMh8oBoYRMLcaDLhWmZ6/
mwU3HdUpfgUsouaSm08VvhbUdcs7ervL5ZUxMVSJ5WaF0Q17JPxfMxD9wW3exIPDaknOktdAeHzm
xvWjKuxNDOG8IHzFfh4mS1wLWCJCabtzN5dp+O5SDlzP1dXn7/sBt/SbeT92LzXUNQ2LdedR8Wnw
QBaUpI4B9E38BF9iWRX42VXH0XHURnK1ggCbkyArYcDj3d4z/8pPg8Qfu7MThMCMwQhCiV6AivzA
nKREHsVrrA938cD5Uvj41u1hxr/G7cJ9NNtSyp1r3sr9dJeOGw8Aav9tLwd7LXf4sbIKQzCM1bUq
KaU4sqgKX6LllcH3C049aJmNapp4efYMJpMy9Ch+HV7dG11DJwzkTw2AOAA+71UUct1bS3hvTR9F
T6chbDS9onnu0Wht5+nUqKC7A8SX+M1HiijiWn4oOFHwO9VB5SJM7HqTUDw95BK2bluluwaC2yW4
dbJgOEG2kBWuPQTfC5BcKk+4m1tacB7QKR73iJljq3py2CkFkoMrdG2pfI+V0u+9eKxS0x+6OXax
jflTIqdDLYFaDdK85gTR0evwfexU+7UPoutuhzI9JgWy/NYblQS1nQGVW4iHKALieE9lGcvWWZYZ
OgFbfCa2prtyRjSyPAzYHDbfoE/2lZTe/AhJ6VctwV3K13SawXcdrpq/MD1yd2zUSRziUh/v9Ko7
UP5M3GgIE1J+Mz+1jt51x1xZzeaydaj7DzNvcVbrynF16Q5jGAjKof6IUFQTCK2uKNQHOFeN3SDp
b3TXBdX/xp4XiXxDNjcolr1XP/Qgy+n6j/yHhuPCPWo/tvMkk0gV32Volum07SfD3sycBJCzcxdn
0irwYx9Dz2ik6ycVUMZZOg0gT10Er3saoF+3cMiivV7vjOXmBdjMuqKxVHXBCNvjmxmRo1LZvQ2S
yaAnUy1u/s2JywNQGpny/wCrVJL+pp/GmK4zHGSSkRNR4b/y7kuh5DVMSXirxV48FVSGMhRxQIlc
HHtkxnlH4m2LVZ7A8xzZBICgxmbXrvLHndjFzIuDJiC1hIPnsA5RkW8J9J451AEHZ/hyVpmjdOTp
kSpngY/CwVRPwIACuhDjNngKMuHWdsH17Ex3ExRENbaxzYXMPxpugi/yHdhTA3uywlMm4R1X9b/T
wYfmc1LUJmhYPj/v/jv3xZKEXeu6OR0ZVqn6aMdoeIiAlpx9vNIHeC0oXaumKmesIU9ZKCbiD6Il
BFU9z28hS03udGEs5uUPRdvSKEmK2aaW4AurUVYcqNGzzbeNM1t2SAlodno7CF+mRQidj5fyv7+d
VzzoPtMoe8W9MI0/8Jdf/RDmgsk+2CovPtHb6sii4LNaEatUm4QLM2801eLcjrVFueVXbNbN0WOT
eO4TMBU1DJ4295zGz3zwOsMQRfmXLNr+lqdaVrlzoZr82WhcQmDKwcUoZ1c29Niwb9MrFw0hhYMw
f4/SVNj1DUPBaneloY1o0HnTc3TAsr8DFl3oJ01i/1YAApiXz8xqm4ps/SHS0F4xkvlwl/on6XTn
xlOGJgqsU3pDh/UInKW1cdSWLV0WIKNBEyMJfbp6lN39qr4BPh8glnfw0g8BowF/A4h3qlWinaih
Bt2HUXmGOw5YCpl9ly963MMowOOkvTxGggI4NtfZ/+qVKZAMd9Q3p7fV0O/wCLhDJl5xhKFtCuhr
C72/jbRDwEKgTwf3CVas4KcrN/ksT9A5InqWC3ZVXx+oKnydvqxt2e3mBjl42aMiiXQNeutqLv1z
Y8yb13/JrToXT7Lh7s+tNhucu9x0ONFfhoJ7RF0fkWA5AoVfeFW8OhwQQcMK2Qir4efP2/vbs7RM
V8V//itgbmVjeX8VSf7IQezoBcPxAJo4AahPJCaLsWjyL8vD9RjvIj+3Pb8GaUPPfQlFw6qq9Gfm
kDaPO3ZyvBUzZnAaAKAhDT1yeCAdDSlQvQCweyrOIzMMniPw/eformNiKWAa+0zhu9XqYAE8LFFz
4GJ3ND8kRbX/rnGbNEDox9SdESUttkRuDubPv0u5Ss5HE2C1f7KeHIRpnaBS8v3KkzZYhnWTLoVm
Bhf4k7cFcQIJ7FIV/fchQXfbjCR8uidow/g6XBmG3YKErpqFR2G7AdSUPVmrdTYS06lXLhqVQylB
kN0zVyN02vxlRzuLJjnJ5sOxatPr9pDhDac9W2CilcV5I62RUzN9HRcO9k7Z9wuYb/U09JntAMea
0RW1skTRCuWHNW6j6Gmw98BAW6m3hAm3ZhT1kAdUcFJHaG1fu3wT73dhSBYkAbsHNVZ5PIvWPVDA
C8JhRnfdJ2jUX4yF1V+1hkIrVCZGkfA6cpCwjRgBppE4VZmyUdt5Nse3G8ZfcODc8h3KsPqhpy6b
bg/QlyxyDcCmMJSqRq4jwXjfFNhw6IzxRrdl/Jps7CpAYsNfHJz79LimBxdfSHESzsNkh65EHWNL
slTYOVWek/UfXRlbs9zv8i9L+ieF8P5+u5iq9EzI6Ku911XuEFd3rFyUyonGDlpfjf5YTITl+MJM
HjPhNhrh3qrFW3Bq72wiFNttNlVcx/u5YPp/ZgEZtQvdxYXek/s+xEwYo/nUlnTB2SXRkz1cTJrP
/ES5Xqdcik7RywpHlcVIzAB4zk7CJaJGWsLgsrp3NnzqxvRJraZFcI/CNp7OcYmZIDCqnI8ssGPP
9asTrxO29Mg9yEJTKxFIR6lmEWFedwlTuUGAnrzrfel/uty2OHCtUlqraLxCPE1SJcRsLKvylmuZ
beM83EXAdMVdif1JJbqcDC9VKkVDEm1a+YWNnp0VFSr/6vwcbKuPX2AI8XsLGKJwfLtbqJ50w30F
VGmuRl4izfCX2vXlH+7/f9FKQLjk6yrWH8u4DF6ekHa9jKeQcguKztS3aTDq3n+Wkqa+CkYFYL2T
P2d+FkzUVwHKG/mnBaqV0lL23Oi0c1FovKRzYZXY2IIR0h+O1wTFPMKiOPNyWgbmkIT4egH2hiji
kSDPC9tpFgCsC3oJY7YyaY/WBxc6y7x8KU0fxiFvDUzj5db/8g2ycST+hnpNPiUQ41Cnj7m0Ogje
rp0mJpeVylVCMfAOc6amEsMMORIM5geK3nOIv4YFF/7F8Z1HqqTpI8vq2GZN+xSA+9UsbxuRiDig
GVnbsbBzreoPv3ljY6LZVbfoSNaSy03QYgt5zp376chR/BKjjj45UJz6P5w3YIuBi/A40n4CaS7x
WTt/4JA9g/m4ETrSEgSxWDBpOnkKP/t+E5vwM9ztfFAXuEuZPSf0GY2yBc0bnr6pCkCHWVV1RLD0
uZi6/BmJpO9m/I8EyRjz4gIq5jsjJDk8u2SOsZnCQojxo5M8sOfdjoemkzfbW667Y5nWPYz3w7si
qk4exqPAocgnqe2c30fBCk+oiQXk5ICb9oYa0fhEyjj/2vpVYhw42xq6MVfkv2A9k7Ub7+KpbGoC
l6F1EkNtjNY5kIomOGw2kOSOuBJmnkx8l/fzX8Iv4xVhDmGKVV/y+aqGJWnmAMY+WyK4SKvuAtkD
JgAK+bcKSG81wPQAkaLvdWl8hLIyvG6R4X+596+FHq1rkRAoPBuwtaCpejFDgDvgfagvNKUq6n0c
5MqxXG4F/zhvQJMDohBHYWcPcwPMblvuYeS3yPP48xBJmiB3Yvbs9lwDYCbmwybvx9D0CBYDbuES
iiSoUongQxMtv84waRfsWVszOdM8cJ+T+BFO11qnYXxygRznObjUr4c4cqlgcQXRm6A+YfUdIakR
4Q3uDFzFbCv4Jl0AY/Q/frYeCyw6TWXHk5WsEnIJ1ODh6zjH/F3AtCp4VjHMWeIUrjB/zAVaO4Ny
MVHz75TT9+ltvmQaC8DM0bbO40ojWb9Thlg6i9cTlq0X5uYCrvocgqKRIisSz6KEKoYWKyJ41p2H
NQGHnnwxGALacmSMf/TVyko7PBJZxUbbQrZlNhAFe9rqj1j47rjDrVsNkumtDfcru1pOUdC/3jzn
XMvSCSZggWlk1qFiCl9cdo0Uun+lblLHiJVSDihvTCsOPh4S5wUNZnUiXD9FN+FvnSCzblRieEq4
7tnkOvNmMjdUIieR6+NY7y1c0xdm38Qp+fLG+r5vJXrj5j4/3qqmkJ57KP6GclbaK9ABOHQ3IDtU
K3uKE5UggiDm4Hlv2BdLy5IdDQXVV9sR0n3mgHIbC8ahrx9dtI0ZrqPsqZaymWU5BWx8Yp44pRcs
90X3MG055JDIMopwKvKHpCEfzFjsoZn+Rq7MlLDLI4tBRvp+pNlI0ApYJUcEI9gyt9n+oKlO8LjB
VfO//JQDeGm0p1Jc5Txjz0mc5Hnv8eX8zXT7EihFn8s+kcGnFdriPmJvfQ5cJAfma5nyx/2rnyPV
TtJ8n8vO21v4cneWBhKb9q6A8bZp2aIzQYdTibPZM3qMTsgJU3pr9kiNcrpcFvLLw2Qq2qFguvO+
trX99qTy1pY1SISYpQ4SxuZuXnSP0VgOD6qv8zHCopYvBlyOgsUnATJPwzUKzcNvDQfa5IQh03Pm
h7X7VCF2cKuriC7/St56KaZc3t+JnXeGeVEBYHOrxuMQ/NR3lp3PezA0+qzlxxCiYhZv/YBHKbuo
BWRfkGaNCPBEmoNMZxCkM7+5yzZKMSFPt+nl88F/4Ig8ePsfmnDWC54Kpo45tETlt0m2818agjwF
pcRWG2TMIM5RbPitIkZDQ3/CNu5bVhIUw7jRxIJ18zMSCKr+VUzmOV2Yfz7WHSIknTaMLW/3ahnx
uAvjtkLcGJ2izv8BpnlQdxkrp1fOcm6TIH3RnqPEOtTt3uclov/hlSwNwT8pR0+Wf3WgoSMFuvP8
RpwIUob2AaLlqSOAYrVi83Ly/86636g22j9/swTVH0xcnEIaGzaVK0m/cazWL9g2pyleDMbgUixW
+ztG15aYiiQF6gqbpx7fs+2b0osgynXOIL4+LKs0wTUfNuUFftds/9eONFYO/MxrrCtodJTdfIFt
U8MHnHZ2n1rSGt+9MAxB8UJT7uUOL800kSumV5Q6G4HCYkbVHzHriXf8em/kAEnwIBoJRwE5Pxm+
y21coYZocvxHj6vjw1V3lQswSeh4dzxwUGr7pxS7MpiDxl2qsT+ut20fwCP1XKJyty2hVO0qKGZa
D/3v1BF4OgDka5pFlmM5+0YXdGI+LoYitFb8eZrwfQ8PfcMOlKXrLho8ulMzF7fbCV/l4w6VdjX9
Rb5b/ug0wpE/rjc9jIwRFfodtiqxVoVJVq5p91I9xsbbq1Skugy0iM/1L4AX8lzS4IPcGeNtdBnq
+v2K0+Hkn0l1yWTV7/IY+02w30+VsMfg8UpE+E4i+CQmlbZ4WeIssH2JA6K3NtMTR2O5+AWCtZbF
HD5iwDqvRVm+12ojcnJ2i5HZhiFt0pCXMDjkxZyJSFHl3QLPBR+4/7JJxDkhvEG2YWZnVvIIqD2h
xogxQrg8rji/clRY/l+l2BiNdlOWc+TCnerE9O7U75hvrr5SuXdNeSEFo/bl8Cm4CkLm9PiZhMnC
cjGEcMK928I9sKH4pmVCzkjTIDyqOpMJBOx2F40rRuvbB/TGoef9Dv7o6RnfrCa0KrFiUYyn1SmV
vY6NflNrg8QcifAZ7FOLfWd4kDRZigLW/o76V7qRRBX9ZV1Tp0JeBK+GK4A+0iZsu0dD3XqsrGCk
pmNFn932HYFkHFaR+oGZdWCaCaIH+9WBfciFZQoUomUdb6tgFdrRtTJB8wnHUhJs3e5g6fsIIPWG
RtUke1LukeCVc//B0E6V55J7jBEZFP+gudPQPu7Ay43nJbEMk8h7F+raIWE8nD3Y6yM4QqlkAnT1
TxKIENqjueAC+43q7uTGfl+40mrnimKZHJ7y873d2f8qlFkWca6I/CSGBxbRT+CQ/wCJRjottq8t
EAnyNOboEIdbQglgTxySR+2aiKJn3V/na5uNbRTVjAXC/eiX3DVbz37urdsio0HicJB+v/3j4Q/v
WjHn/bPgZDmUWdp093+i9unrqRD1kqQgJkpyZE2sBis+50qlt97ZeKO/TCu+1YqzU05mE6GEYZ3J
nHXYM8LxxqVDFb8bIOJ0llOCiV22IG/ahG2zl8/UX13t1MTHMqndTvi2bSwcTs08GqLouR0jPOqh
JuaZ424tCABYJjYmrAUlXdccwEicb8P8ONutg8x3IBbU/KDxuWjtDiQjSHRfXQ1HbmYwuYG8C4rK
G1ZosJjWOz6R8yv3DfWf2q91qBnFiYwFUHiODSmgBec5HXn6Zt5datby28qynsXyrNk9xnto948+
DFXffkOtxNYWqz4vG0/37bvCcqinX4WLuEtxuNSws31aqcPdWAt7vEylArZoliNKnmrjhwt53vRs
etZ2wNiErqRPjXsoexLAFXFlJ0t8Qu1ymr8ktns+lurQrxtv10GfKQykl6xmBV7g/5FeR173d+ad
EMGJAN+QRs4oyNz5c0TRCVCiIW6d46WVGuDDB+Pagu4QjxjHv9nA6tAlf0AVdAxqwrP/dN2Ivhxf
kEKJxpd5RHGd71jdZocViS192EzmLsGjvEekA+T1TxYN/cICu6ikEA9kWAAaXm7GpZLuylyXfqed
VfcOQ5j3jFoLDCyoonnz+N51Z69rBpigEUv+AcKskNhWREntopcKMvhATXZzXhBcL3m9zoZ7aUVi
FyryOdUunnrTUaAV60c9UU7Q+8tXzAyEejYBmdiV7xdHDdBVDmJN1f5fPSxTKpHC4nm/9oNi9GQJ
ivTj4AmtIgoGbjk08ZeXqnqzsYk2ucvKNS7SWbPeYjuScpO31vq7i1CJ9NMijjGgYdCo+YinrRc7
OSqCEimxMMD3psEJw4H3w1U8kuBmqXKt108Cw3zpKu7uNIe6pg+xGYo6x7HfbxnI5KsfjwsVIEkO
p19a5+awCRPnTaYzUArU9Lqc77ddY6xjTqTBofvf45IEeoB1233DijlAUc+MdEQO6OWNfMtwEfFd
7RCiwx4aCz8EPAOC0hAtV40/v1H3tms1EoiY6V6CxTdU4WGaNuj/8OcSkmYr1q5ewvKYjPoCt7ek
R4Sf9zc92Cp3c9gJcoV3+Fw1dq62F1l/GmBNg0utKPWQH2ahaaLjX+QwbxhxXG6YNR3eQuHLUEFF
AJKo9wACBSN5TyUvMIPROvBmElB2gOhhP0FfXgrmkKlxQZvn8HBuHyOVRIg9SBo3DM+1Ux8tftTC
rFhRb2I4jYf8dejvW7L4fsHCbzBrDsG9N6x2gLb0k1RNiydHifA5odK9rCcEPhT6o5PVgAPDwozK
eJcif8JGoizq6syHyTvydEH3Gwd9zm3emb9CnY1Wuj5xkd6bkGhhEUOHuQJY7aLNvJRz1FUzlY8U
33J1S63c4E/fEZXd2jp3abIDe9a1JNDkKV4ezEByw67NNwi6zhrasyIqfDa3rsfSN1O11YJDWxI2
dl+0iVVdOCoLIjkHCJw3wcxo4Q3pMh3Rc5t8xYksnXdD9MFV6bB0HDh8iUT+24KOeD1nNQLeTVoq
cOzllF7lNGanRRGU+1T372QORpdTOKDW9L5X7CJof2q2uHJPmx4ZGLvVqzWNXormUYv4QbTaq1RG
Mcvft6hApKtnsS8W6wJB4rKL61JkmnSl/w/uq0kLiKo7AFVDtOCUFkYC1IS5LHVrNhhwiK7+6ejC
Kibi43Wmw9ZYsRlCrp1W95ERh4e/JiN+5ak577wHu5KRXD2Y0j/eeDRbJRj2rrOOdb/USwWxvtLE
bYQdO2TPEAvDwW9fGf5EPiC8TMckPj4B4T/qxlOGFp7HS7O9kwtjPjhrxatGkqmHQ9S1IGRsKdsa
02IkbqoeQVmqZIbvgjszz2pVo45olv65hJLgkDjDad7sqr/QwOwOBSwTzIishSElidCFTH6zYB+b
6EczTOcURxKoPpspolQjZ9Ok5zFHuL6sCUdq0sG09BccOlyVxuMiIC139dXWd5O5SUM/mHo246ap
uxbpNXYezBErTMiGO4PAH5sZ99Zcu/xBdCxoQy35Uc5VT270QlJfhds4y5pv6eUFp/d5kokdTjiT
JeTjjuPQa2m95s+K+0SOxOV6BaJuTDn6nkiwufJN7ASGT9F0ooLQFuzFn80BrxlH/T99KIlkRnig
Jkrj46Ac26UjWKVmbi2niJ6g1bMv7UrXO2KqALDVI0ufA8B/0NHNhxL/J/EaA+p4DkVwTdECT//h
roogwVce8QVxr3sJrpMGXXfU5GglirRrT58dAq94FgoaJibn2Bs2Tsis0HlZUXdnBUPnBds7jU+Z
O3zIOH+z9Bs9xwS91IfboygbrabIOMQWaYpK+PZeLLC4ODe4ThyaC3ZvXByMkeDTf8aVAl8im21o
ledcofYPfxAdOUvLvpYVnJM9tKPM6acyYGQ7p3EC+awOEFJIG0Uet9ZePrtsiviYjRCEs/m0NSv2
oCz1JBi5Agcx+8qp0fQvpSJ70mdwjHQQBIYiTkd3pYZF68c8oYDDqQrSFqhDDUZv2TYmZ8MnPyw8
7/aq7Z+4PDPOyk9IPQgXOn7u9+hzq8SEq8EEOX0+WvF+SPqxWSKJOpk/GVAvepywUkAwIWf7ogCw
1kzAAx19rwRHSUSotTtmXyw01VPP35vgJNGKhIGYsQeidu7myJXJu3+aRsiGgToWO3XnZ8C3QnPN
hpUZAdUmfEnveh2OE8YyjymXGjulcsgKnQZS+R9d6pHBMuq/8sCJkeLbYER0Kfywj3xe5uSQEFi4
0oPWdookGtbqohszHS3Ag0tcPytxklsfzxOq6wIsQb12ANRj0eoF+tSJaPTHQaYiJzDUwVJn35Gr
6rPwGxPIpJo1Kv172rj6kP/8vig63kFdKcujvD0eLVSIh4LBRAh98XDfA1NvlzbiFYiYk7MDNyus
IWLsXOwIxaHjCXiRKlM232cxwuBFNe6m8llgJe2oq50tsjW+uupiDksFeJ3n3IdUOzqKUK0Lvc9C
ej3puG9bOK6tCTdPgKyq7baiazVLFzRZ/4jpjxf7sqqhGP8BQkswRQwV0AydOWXI1MXDVsj2/qLp
RWpElyySgiuIplmAMwg37oPnubA7SEn9UwdEkO30+1fCbuUCoeHkCcZLp68KhdLTjhg4o9bnnkwK
JcSZZqLIj4wr5HtwX+iajB4tlvY1hs6HQU19AM+9WcsR0EM/Bp7i3UjIZeJwjmKklaNq1lNREBLv
hKWcQW2WZvj9/Yg7W6mwmoRQ6TNV0FRYt54vdEbgqyLe2x0EnPP4YkIgNC5NYTylVn5J7jgYt+Cr
n5plJP+TlhpD4Q0W8dSbjKg/i76icW2xBCqzeo7Z8jrJ9pJ4L+Iznx1fgbyjgWhtwCjkPWk415JT
cnJ3r2pezrG96Iw2TtXnSfBfVvVzk6+F0KvVNxwpfpfWmrPDXR0qwXhK3MLD3rKt8Gls4Z+wl/4i
AOWMSGQOXX4XWel5WMywqUL1YRe0U1NykGsrOmTeYU/hPhCDyC+zORMI2kh5losq4fB9OYem8nb5
Xs/FKQybHQ1B9k4Xv201ZAoFB1YQz4PAF5F29V6CDy6/cfr3+BoyNVJwNO72DVFW1a5oPoea9vPI
34QGKn0e78VDXlpZ9wA1W+Bca7+IN/hHaiBtZN0WtXUePxeWAozBEf3EuOSdDlseM0bnRHECThJU
CgydJDmc4VYHLS2KyUNPKmf6YsbNxfjZarOWzajNai8xQ/GPFjrBFXuF1fXFWsew661QvLpHLFfa
WLN29aBJat9KHOE6nI+15dXjCCNKpSBmzaE8PI967PTK5fGHolFICDod5lzaRJ3cf/n2nFkWVl14
/u4lJYhLD4HNPzNXVqouxBT5ZwQKZJMU/1dfV3aE/KiG1zFtOWWy/zSWw44axqzLRhIB9+NTBoZR
jRkKhkqBH1vlccMM+ic+VD8+CqP8OhsMlI3xtZ1oDjmJaO8v0FOyy0vqzrJ0dB9Rs2WkhjSLGEUa
MaWdUKMG9BL7axgTvjVatTPfNvViDzpGoDjRmQSJwuUseAybvWCOsukLIiQA0WVXoy2BF4K/tthu
2PFP4bCQWpb4ySU7f9Awdz5ukTGot167akGH2/Dc9fbn8S244AHlzh2xifnVZfuEMh19EYImZduG
pbq51R+FfyhuJEFO3TUGZapRgQlljca3S91iw377PtYfBqUGhFgFWSNE70zFlBS2Hh+hrEYBjdPn
l/k47cwktgHatb3jz+m/b5S5ysN/JHcc8jxmLZ6A7tMM68DB9ULHyjYwI/fGIOA94G8YW4UoygAW
WzLDrwPUZ4k+fSpTnTNyAZ07O6HC9pAVJPCS9F2G1PFsrQHZLWG6WsiaJ+qZOv1Pw5qnD8aIc6qs
8Mezdx5Zb+DnzUfamu8qOCvuP3RpxyNGoOnmQ52Btf8LT/gIqXrwU6dsJYwwiI/AWTjEHA8HHN8H
M0xixtt/XPDmJkcEANvdsclpE4PffwMeZW3L+AV7tGGXmBf5QfokWfk97iHMxOdIn8ORvV30IfaW
EpBJyGbnY1+aj2cYEcJuyFd8ZE5EkxhYj7eX/DItA/onPcl6FQ9wdRCoUM7uyDZhD27PxJT13NAm
47iycTCbnJ+Z1OD/CiZHv49+hjWsffGYIbbHYBXhynM3Jg2h8/K9JL/d7AFZdAgRIGV2aHFEgkBU
cxv8pIILjAGomvJuCPi17TPMc+CA+eF/Bo47gcXzx5/rUy6z1KXGhPtAuCmq+F0GdTaFG50KhYKF
za6VTMtzp9VSA8jDufTuxoe11d7g8X5LNwI53IzW0oItTUHdQqRivaMXf2ynQV2RU2el/JF8FsLP
EbOkPZB11stNBbFl95fg1cAobjqJ1fg/KbQE3KhqLJNh2xPxFDKXcxss2mHZaagn4s/Be25FDAAv
N43wyr+UK4q6dPiZu8iD/XlJRGFE2XIQe4NjKSTHbWemeaJEKx6DpmneFeaYkYrkewG8fGy5vy7Y
jps9Ar2JMzgTncLWTzLEDeZKZB8FyLI4sSBrHbELGUs8lwpf4OgHfJCqhLaFw33RWCD95U8lq2eD
r0stzsxBOR+I0NlYQkr6rerJwTFwgfOS7WfFdz3V6wmCcUdNbL7xoof7ekduiy6cPv88rMurRQEu
unkDyaPatL8y4ycKuycNT//eFlFamulNr8pXyUT3UzJykEt+23Tq1qXGQPpViNvXAUWYRBarQ9/S
vqc3ml0n/XvQrX1ysswB+vEkJF4Qf44Tsd1kOY7BSOUrOZ2472jTCDkt7Pw/yki1qggL8Y+eefHB
ZorI+fyEghT7FmCubXUQGyd+95PwwTHSzwVLn/sXPu9cwRD3HB+c5Y4n3ZXVUdp1b8klDRvCFup9
bWl5NId12isp0ziL/kkC7KTSpcBdmkHmGsewMbdV83k5Alb7/G39GAPvo2+kOP11dVGYIQtsx45u
OoIyc4udc9Qmfhv2KOY4jZCCc22Db+48ViA1K9ykxCri3hqC7HVFkrGq/XvvFFi4VvzxRK9rLg1f
J6lDlUwbl+tPQz6l1AoRZ0m60j43eB8D1jENfgIjMbxKfX1iS556wYQn2UmQVvi5fch/0GsFw+18
OTf2cdG9xEQ6Jx8rToeEzW8DeuZWkasNBAv25eW1jNW0/VKw1sfES+ke07QXOO+Vv7IHzUbRf2er
BvSKnqfCQTDl9zHaGOb5UE1NIo79lpYQ7DpUxJOLLD0Rlr3PaGbB/ia4xhtBd3c+4o6XdGAEH5Ef
EIK3MztQd42q0b+av8oOmby+XKPPhnvuITjL+waus0Mwy100eSgKt9blBPg5g700nzIr0eRNX0Sk
HemWgrDChr1rcPpYWgmszN/6/J+u/0vWe/EyVWIgDeaTT+2l4WXgIE4NAsq+gcowkjcR30FY2Vlq
rlLWUsqp43fLDfFIVPwAc/SofPvjKH0Fi7rHKH29o53FnejEjOZMWP+nS0tVNNbGhZPVz2y8IwPN
5An96wFURFmZl1Elghxo5Aa7pSs2ls8EkWgT2NZdQP2ZwaYYij8U+ewH2ZSYQhmoHlEb76sUp4FC
cj6y201Mpncn5xvojlOKmRdiMS1vsLhgdRu5rX+Ax8XanU/Zdaz82oH1Jb6HAxBsnrb09wC8puIL
j/XedauiW5yeHiHc4327d8o9dxD4pGzlvCFSvObKdvMOf45jMZHXpDHLFR6FZ+nW0XjAvgolN0HJ
KQrnnKxTPTjm+Ea0XY0v9D15nnhqxvxsaPSLdhdRwJMH7MkedBDlYjzq7LUxkxYa/rlAEAhvdls/
dx28sXTtZ13D1Xy/9R1BEVcrKK7O7ZjdywPnLMByCu+TK1nBaNzL1djk/2DTFK7CdYya/jznlWQX
uzf2SToOY+e7TqaCWzEZdX59I1peUugGEPOZy5YrNHViBi24tJtj7ATsMrR2G2Qq/sVS8dD+6WKs
Zvm8RF/6rl4foX0xnwFMXPtQDXeLUvKapyYb+7+4EEX9XXDDHfPap+wEQruICsdwPyq4OoNQO1oq
+BdsTQ2ag89NOQoD8Pu/9ZiXf+o0aWHlOkXhuTy58h6vW0Soyi6LKl6eHo9aN0W2HDxdTC442msC
gqgMGwQzC71ir7NEhfb0qGY3tcEwnKJHJjzsbZMIBFg3AjtScF0pGXcMLWSEFaP9wnLWcX2s/SIZ
nkus/plCDnISYr9p7t9hgTCQqmR1HK8yTDVuHag2GQrq3dfQVt747OBn/iGqzfP6VohuSEwQZHmb
na28FwM8FseZpcqFaMPi+Xqe1Z/mmAQNfSCi+vlsXNGZMLBRjvlsEJOb9vyt2jN7qxGv77IvVKaj
sclEtOqFg+3H8OlI7pGFC9MEdxe37nvEkN1v+UaZDQErXq3QLRseYI/omnDNVy/Q1SC2tvTAPGuR
IQ/xCPypFfpo5dkd3aoqZ24olN14uJvkUo+w2tcetPjZGYtR0AviXGIqbYvkY7zAWPpE3UIfqaKZ
VM+u+/aCEAOQEx90Li4Ix3TXUEqEaVHOAWL5POGuC1imfBUHv5aLCl730YJP8Bw7Jr6M9mvhNkhT
Al9HUZF/2hEh8+NJidenN8PB8DscWsfIoL7sVFnN1hWI5nadv7/1HqDigswK9tTVFnBDVZkK37HY
N7G+Dhvdyn0z+WvN56VuqLXqpkoFk3wuYKKVQY55jaGlupestBMW/BDVXgf2xli7sX6LzZaWZaBE
d/MjE+zIHT/RNpIbVNkI9IE1tiG9F3eLJ0JBifa9sKHffa9j5paWZUSdVv7RmxNOGArxkG/u75yn
7BJ/tWRNoTACTTpraiN4W6wNCriBnG9JkJ+b9esOzDrfn+5y+y3UDflrA8wUE16DUlD4WI+oavnu
CuEfhFG9QypZfWIh7h1L9DmPsnBIuT0bTZTHUiGTjw9LDDrSzCvD+EFQdDCs9r6UHd1lNZL58TkD
/Bkm/nsDPEu6AQmzsen4Lc5x1g/xnV34sTP3PY3KLp170VHNYHu4KtntzJDVdm2jLMygkv2B+N32
eYXErKWE0+DUEGn8rc20w8xHQgRPQwLUsFFf0PZvGTI+Zq1U4qYeeb+f34bKvijHMeE+NfHheNMS
pyC8nEvb+O04Bp1vJ3COzGQnI5jySIaWQKiLEbXyaH5IiitKzTU+di94V0S2ls3qgsmxa5G7l7bL
Xl0JUqv2zuzBMsv3FYOsqOPNrSvlQN2LJawrAbvLOn7EpdA8sIv3Ty/P+0+dKm87FEaaTUt3cNZR
iKZX2CbzocmOWjJjcRhYeFJfohBWiyoKCIHhm729vSDMVuTO9aVh9EXKgjqQ8jC3N6mfqTs1qfL6
s9yQMdRuBkoFVdrTrYJ/CYawASiLpsyHQ27CyMsATXwRmUot5k7NxAWZn3ggS5Kv0e5oyDy/jjx7
hggrMDI1CoVkOl4hjwBTDnjGAMRrzs9DBgwoK7shHTiRp7SS1KxzwDbIso/hrB4FF9iuK6vt2TGF
gOoyBvVXoLG0tJvw/eD0ZKJ1J6msNJtS4yyrSuBo2QHClVHad+9KcdzQWffTV6Xs9JQV7klXiubv
ZQa+6U5brYuzUXZxFF7/iqusxAbtCGAbkE4LoZtFfHSeLv3hMosqr5Vs97f191SEaxcPymeFx8Dk
6JDbPeBZmjAbolsxKGODMKJjK/kdtN6FZlFpfvqNyZsDghQ31LEcz8pzFmqN7iNKuMCwUYFBn+0l
ANwYtqOEipmOBAC+yT94J32KQm/grtW0t1FUXmWECuUci6OP8CjMqdSr6V5HnjfSRvMgmNupLT/f
C+JOkLnl8M/ULb+yd9ZYP+h1nWEDMYmapgB8r+uwOQaXuTQK1eBGFUBl3/54UxoVBg01kfEVWMm+
Pq1hJLfmeEk15lMqLw9Y0CQdYO82sPAGStm0sJ4i72ElhaSWtez2x9fe53wIAT6ogShODEMh8ADP
avBiQjiKTWljWHT22CjDTegOB+7yZoUAEvbIVt7RwIZG70yXdAvQnZUkxULQkKcXtowihLSiFYej
8aElLGQeNqD7ADsK3ng643h4uX7WdpDZBvBlgpxoCBorRRwwmmVpXkwvPwB+a1gReTJ2Zf452Q64
0m+qFjJrLV5Pb7pSc8RGt167RG5rtcOAsOMO3bwjHvl2DztUj0z6mVWOxl6B5esEhlghYrLNH3ib
958sZls61BiWBKmJJK4wo//m+6uHDryADNIpR6P2zYo2LcqE7C+GK9j0pyfQI9tf3mbPn055PoyJ
BeHbJib8ifmm4QlO/XCAvMe+12bkYqsEIJnz0WLYVDjgAsiuGHNKWtCmy29MOBV7F9mEHCg2NPKv
07Rxv6qwR1HFaI/9VPGtwndTli5igI4N5pAD6yF3uuXvtrMKuuHp9Cop8AIHwHXHKg4dnh2qDSYK
XLJok1v66YohGc1Jo61DKRcZ7Yg+rOEjvmLqSl/aJw5Op+GTDDBX1kLul2mPBv0gu162tkJnX1Nr
aLS10Bf0JJWsA6boyCI2Ky0N1QI5yN9HbRbqtMvJEZKv9HloKZHVGAmMOXiz3TrLof/aVAYpQJSb
eyMmK0mJdwRKpsJzRafibMPcI4RBUO2GsltZygCCp65yghGHuhcjEw6awsU+N38AURER0PD9Wu28
t3YPiKLsykssJ4CyRbOSYmdAWTwzmvvM3QT3T0MApoLo55O+sdXttip/WHr4vAFT8eYMUmA9JGyo
QTsXHNx4bUWeqS9G181cW8W4DHM9IBVF6Tup+XDOFx4em5TYWcT+OOiT96pRlRVcXxR4SDuwSrdN
zNhqo7VymQ3WwgN1sgycvA7mOMZmgZbqP+ypHN/7b5XYlan1JGOcNv1uCpNH7K3LEzDZ8gTHoRmX
hFky8ENeTBJFSReU3LKnPAD39Q8V7ewJ4tyGwk8TdYWfNWc/E4FM2Bc5g95k042mO7m7HXNnErvs
9mWxK+iH9+NH5HG2p0nVuZCIJVtJ5YK1jPusxnm1UI+JEsOLM1as1NgZUslM4t+z9oZZpnu2FlRB
ZA7i1/Dk0e20rfyxecTB4TiKQNE0EikQgHrBYAL/UghLow5LA/CvSItLB7ZhDuCJN0lUwT+xLDQD
epzvD8uR75Z6NVLFRHIUOcZK1w0vzDtw/I13d7jG03Y9KaxA/i83Cs9Nzc0jhb/o+4/30RM0zlYZ
DcLsuyApfXyxs52TIGD6mb9gaMm3wKgIz2jM6umjyy8z08HSD42xboOJwGUk/Ta3p62VA3rpQAdg
LseD5tPyPjU86s2Q/sdQpWO3eY8uqnoqHyxHXEFHOPdfU/pB1gXcLFuQ96tuQUn0KimXur5Ox87R
ovlsEPky0ICGvGy2cwj4BMeAv6h6tyPdMwTcB4xdgPyib9NSr01Yd+rSluy1Snk6ktVsVIY/nz3E
y9Ugqjhp+/4205rVgdLeOoU2z7vEmsds4YCJTkicnKJqP2IpWAKYmSlEJmdyUrRfdtANKGPSYvJK
6nrLGNjCk+HakYTLyQNFfW7eV0LmVGoZQprj8OIpT2g1uq/o0mamlJ3nkQEPIuiSgDdL1BR39o+V
s4+ulb3mknO1pngksVTuHBMN11oy0cEweB65Tef3OpDDi9VOauR1DCOIfYP3CF864CgBF0/cY55I
G9M8ms0R5XB6P4Y4SvJFO99qCcr8pbmRpX1FpwtVc0PhX7U03NiqtG/+QfCxjLahKmnPyEe38oHc
yIFskuUjUsJxamosYZ0jZnf7E44w0SJ6GzMJInFnhQW6RT95exsNRnMyx+VP2cojw3K/EhzgYL49
ipFws+paJ0o+i672GpaiZhjNSW9bxXgUGfuh60/LiC+JkWv9tmFlZ+q9VcS04fmRrFVgQElyvJPe
Y8hXO4bQRIqCutKkRttn7fsJNCJIP3nDdxXf+f9CD9T27PxFMHFLcpIY1Arohn8gXCe/0K9tz21V
l4dkmn4iniv7gMjDgwU9Gu+4k5vWy4vJPVKzvZCHUbC4ebHYTfj0TlSpRnFYm5cWFyI2tjSKF7DO
Qaw+j/KKNJtRipf8bSrTOpxFQJTJgbjec43j409kWrghrcreF4U7AT0UZB/knLfqunMhPSl5RVLH
60Nc1XDlfxyqlGTekov94I1tczoEbyhW8WPwylmSb84ZWPqDbCPHUPkgb673Podl/qw1s6ToolKn
GGXsjHOCAMgSwCIanavvtkKb58HPdpSbIBdKVdXdMpBYty7jBPdgDG2YHlAuY027OxiOQEbGtuva
ce2l48xiymNNW/EbLDjgWkjqkz6aVAG0Yw2mLVlYl0ZCgKhBv62sfTmHSGEJI+cPI9txZmmjuGC0
OKyPrhOmspwHeSo5fcBC0kRZH8PdzBKlbR3ZDqd9tCyG96A2NpCtr1QsvJE/oC0aVgRjuXmwZYzY
I+nA7LVCbKc6uBKTHW8ZObprO9fpxpgM1mKG7Q77IvmU1x4disocFOlkEAB/4NxBVQ/HxyMZ/L/v
ky4h6dSGORLfKMt8O6ovpwMl2DoIZ8Rqlue8sg4vjDbs7vXjj8BaukZeMv516GDvyjQ2ksugME1n
XEXRxUzEyRRhqW/YnjHn94XBfC3CMSzazOmG0aGibRLmc/mCxwLJ1YlGIEO+B1VCsgd8iJ8AoUZ2
WGlZvli+K4lH+vcckzmwya0peOjtc7SsQ/NHbh8yUYPfiSysDP86LCAI00aPtYEw8d4E96AC0fqT
euRQ02mvDslEz7CUZzfVLsXy3Xtb6YB4hm/Hie5Jn8dnnFu6nF0nzjzU762uzqAcXUKhrXgpR3eh
r0ffuoTFOHZoOS11sh+jHRpZWg7p0nt7KqttsiXRosgk+DgpqEwftCFxX5ffkZiCjiWx5oNWEWaX
K6lhIRf3Xoq4Q/xJ13cMFYpOOCpjfacdp+hLsfQS2PYloNg5s2P//qtjlhQjVKvfsKzHvVQG81uU
/0df1FVrdapzlGD6rb9TQmO6j2oQFturAJPtSm5lDTmgxil2WmSqD1X2F6a+jzQxl2xVJ3FFL2TF
UDUueNrUxn/Z7CRdtj3t1tVlsetu4LhpicFaE6bJpucR5lPm0TW2gn/eB1+5homPJwCDOP0AOMdQ
MNmiw+kgWecjpKGUr2HFCDBU8XaOgnxMhRou0UxaR9ly8L6KmR4hf02gaQrz/Be+yGt5yGU2gtHx
/7NOVvHlowWN8rO6i6qcAVtwe3DHLM/4Y1C8l3t0+AHcT4q5kD+5sxm/Tvu/ljtNIznCKUrJNkJJ
4uWfa882E9kVbTFKUjvfsrHEM99utv+sQAa6HRP1L4mrdUjrNar6OIWefkRCZa7X/MuEeHY486KI
fs+K5724nuMgKtuQ1lkhD6Dq2WkuswJUxHCIVDC5dsu2bXJev4CqjN/PMZvIzDk2AjpXi9n10dpk
e9I5NkI7+sxdSXAZu7sPYMp/eQY7X0e8nDoDv6RTIJHHwOb/pNNmlzdzLGZmBkFh7sBT7ZRD9Cqv
eKt5AGOG0WeOCloP0VkB/UTabwrDBLG4wfzPPURFJSMIshY7EBfDIVImEnGKdyTQBJlqwfc9cHmJ
v2IRP14eHuvg2MVldITipQeZxJ4+XwjF+nDvwNqi8OZFEst1MoBaad3/u9YHcPKxvqNabx0TZrzL
lqAcbAKnq1t3ZB/wnFTyFbefh0IUY0IBwSt/1XfFGZq9g9uCf0iNocb5uYS1apuVw3G4rQ50yDba
3mvaB2PBJIquEwNMcTMOksL2RjdR5/mcEtx/PkaXz/x2U9gFQ5N4uKhJcLsSygaB04XKYXYMrm4U
LQ5rLACkHrhuAr/ZFb+3fJmB+RbbKifASsrZnHIwlp4zL6CKFJtM336Cit1dny6EstSTFLltWZse
lIXQTbDidDEFrBHOKVgC5QpDTnKwi2wUhdPeDjg/fjY2G6ifD66Bg05UNbqKSO1UGLhPJ3U+1NCL
XWRg+a4YYCqADBgiHyTv5C87tXpaLmqF+nOund+VkiaeluQM62HnPo0TZkHu2crlVf9NESqsnbAw
Yc1F3q13T6Rvy1/aDK+u6KzOSnUVink7QctfWLnMON2LDbBwML01dGxQ/SsJnkzl/EOb9Nln3eD9
nvyMrBodVo1mYIkdybOhMudkafu1v0PNll9FnCrHnuUB+eYAv19p3TscsRdC5DZi/OI3oR1GxsTv
1DE1JkTWa1eyG3u7LZJ6C/MR99MgO+6BCYd9p6RcAbYHXpLlB90WLfghDfklHAKyIzLgyM2BqYAd
7wdY6nlatP2Gwm1ynE5acXCabbHSJznlbcew94d6m0Lh0Q61nXayzeGbqiFClIE5XKLLxBApXtBp
ZHpS7yG3etJUXxlDhrW0p94pNcxsXTZhltmnVSsE4ub6Z+4eQf0lnZW+QA/rTRH5aygmAorLMetc
7YA7TzlgsbRQPXhv8t9Hf+3bmFIgnotKE25A1PP/NqYiqf+ROjgHp8yWFXffvy7QVYRFxxhUcYtB
ygS/Ebr0HrZB5GLbPu10urIgIIkQiAlDN+2vuGB1W8T88B7TY7HwZ1fH6g3j18IG5Kw12td2kIzm
l9MgJPlEwaiqC6lCPy2Bd3qzalE8W+M9JHUTsA/1QPZ7qIBwG1HYPrTcTahbBtmuuL97W8MP+VD2
oogRwwZtkF8mcZkQj0+EyZQYMpxCOE37MMG3vW75MrDKfGaGjLeN/VUm3jdRAhDckzfpXV9l31pA
/8/IkzkDZZnKoQ+fSFU626j4+5z7bcxeCAcX21/b0pq2JpstGQ4X5p1M4LJxV5AyC+tCHNyId2p7
/NV1td+D6xaBAR+ZV9f2T8EwqvwJS45A44tPrUoTw8SU/7Jtj6QK1hrmudikPbEhbnPINNUFF+Sb
rh4VkxYCLePOw0cvyjoIvdcuOn8xiVt6P6pAnDHKyL7JER4+8nIu9QiX37/n3m+umTyd+3un2Mug
/dxmvpEmAR2xEOtQdiVoeirM6r4tNDu7WZwte5nknjJr0ZPT3rkiAtRIcu5F7plCf8Wp9TG4dojv
f8uHQUhLE3vEoDWhRAQEtHV2LMq//b3AAqg/Cw7HsBV9UHFl0O+ZWtXRDEKxrkbHBaeiyIiSHhrK
oImwieGwgsjBSmD9MUZcJFOkZiGnuSVDe7eE8bsiHY+SbmiMwhCtlZ10fXeIV1fxoE7zBB2sDgh3
zRcGQlw5tgyYOch1vZrDcij11I/+yFOVO1wy08Ym2lnIeo2QLUH8pL/o5EfbPOs7gjcIDw6OYEDi
KjGlphL1P5izuYnGL1EveMre+uKfab6XqoklgVhg4thGH6kGDXyvT9f4IwWV1IWnM9QLw/0KUzbU
GMQUU6BtWJBkY7NyBSV5nnQghsGr69z8q6Iaz3V67pax6vCZY/Bx62USH84EPSuu4IiVrvr0f24F
uEpEPt8m6zPFizvTJNZdopXWPa07IH9qDohxFyS882nE8gLMhKC0KIW1Y0r8iOS+hPWRQsQvyjFa
8LQfycth6kgJOUNFW4rdy+XsOSYdIZBmyvIiRkOGqoAX5TL3vzL/uWV/bTWhBVh/E6c2TlvhsBwA
YmV1cuMLerBmO8W65h5PPq6Fh/HD52QykfwNR4G7/hxonS0Uau18jyzGIadguzMmHIN6H4MRF+mf
bhSLvgaUp8Mui9jma5zfbmnjq94X3f8gQOeFfJ0emmVQww84AXVOvSyJjkICpbZctbtoml0aJp5w
IT7yqHV1WmfTFqzXGKr6TrYDxPqokdY+s32kKDqX6+m31i+ML1Sa2uiGbVkkJM/yMkP9c9t99uBJ
gVdeHdbnIT7bZp3a4s7yJ5IdiILZSUqqVgBsJDW+SMHYgAPZ+ER/+Ju96CeMPDhafrogW0HKv+sS
odn+cTieedd8BHbmrO9lUY+wKGA434vBD0FPltjINXMb77Sew3LRlLZs8YWxVP6rc/mAoXN32VhA
2MMduaoxSzbcBXjwL03GttQdGU38GQI/gUxCjfcakEouk5Zeo6Po7nUfNaVh2O+5mXAoW7rKJHcU
e02AWxfbTPtFGuxRKeiZr3FRazVTGxfi+n4MRu9CrWWJxWwjtfBuwHc84NMJ6a84pH20A5dNural
5ZKvLIcF6uHiQBCnGLMiMpvAKy58z06L7ZfDctVqvoObaBh3EA6LGWFT0E3U8qQ2I8F7Zf+C/jLy
p9PTvgc6gZoCH3UIzWXo5UULWgx6eo2g74L2MQU4IfqTdhPrpY3US1L6nGPZ23E7XVvjPAjS7dIf
+oGypfRi1/I8mqAyz8XltqgKyR5YclpzKnBEK1h2W5SwFQIarfo35GI5kKQ2E/IFajaryUl/PJT6
EUgxG8DsLFN8ig04VK3U5SJTanL/2jNG0jt2GjSbXgCdTjvarMUioGz6S65mV2MAan9X9xG22KTU
l9kVGjAgIRHss/HJD0b5r3eUO96TWMU4ULYxLaNG3bJEVQ+tOzA6tNtFlltK4rsXMM3J7Ault5oC
bs9lF7op4T0e25seNl09/YjONvxPgIYQzZ1coeT7olS6VhxClS9EKa8GJlLutvS6+Hg6KE6Tjscz
iZB8ulnNGw/nO2c19/VA/gXJWuB5p+mzwiper/vmYWAz1uM0L+yFu3zokYRxQDXMIbYAA1cPExey
LbNXY8BH3I3eduCwGwfUPvI64bxK0OmIiiJQT9ndoykCjgtJyV3srHFDcY5ziyO72w7n5Q3Rytao
yMd4wPCwL4T8omgrVdvh+d4mH/lGhLhNcdsQIsxkcB0II5wcBtdVMmhJntglb33k1Y0RiuO6wccq
xHPhiRgLGn8woE6T39XDZjGVY/b/8gjRRMgqSQpFfPQJNExGXcN9wP6FrjtPvVR28nStmaVkVYOA
vwD8720iwxjMf1f+WkEpe0VvDorrjJ64hOgiloiicDwXZkq+Ypw1qk0utYXunttrl+VX0J9Wqsz+
MdFvUpbu4SrB9AJV3uwVB3lkQPS67FHwC+Y8kcTAc4hcowEjzmnHqkwtCZN1FiegvMlzFTzLio3m
nO1iqUY0gi6HeWF7omSEjBv/eLVYH2qSRMEwLJmOC2PTYSBsQjI7GW0v+7XEww3mV6FaekjNlCN5
yV1wQTN6DY5PqF5WzASLTpIH58ydVsXzsagHoYi7mZ+Qlet+Ec1sX/jZUJuF+uoyPYcojArgUFN6
IvoniL7B/0w3fFYU6uHlEdI7dP+L3rNE0X0oQ/UEy0dRajmD+7fss6DCUvNRpGP2DV5l0D4hA+5B
bZ7psaqcKuHssJRt8fNxEpdiKaWPVLh5PFbCcAJ4XsD9PSAc14bxT8IwBtE+Yp2wt63mXSG7sZrV
bIVVs4pXevSsO7YTXDvohUAMcqzvjN4Twbjz7tDmpZNUVmRc5/CGLGNnivryDcHfV0j4aX1H6HVd
AdSywIm2IBgln7FsxtorkoBPS8zzUU+Cf8RejSg+tPscy5sgego0dk6MNJh2VUSlx2CrQ/Cd45d4
JwwPE59A4Jp/KUa9Z+GpkSy84zBCtx2kVlJ9tDK79Duz7v9W5skU5dDcuDiRg+Olz8GViizOSxuV
NbKcpAsnrd+IxlGa49yjS/OW9LOLvbdXWE44leYmpyiCjMmoIyeK3o52JK5f9MymIw7TXAWJCxgg
E/A88iZMB07jOxq1xv+pkpfhzsRdGUe/dVG4GxKd9WRSBll/qon+E4/a8Uq0wepJrw4jCzFUL7Lx
gF1np7Hdjaj627SWsabtWr+cmIEW81lLZUM1jeOKjqdtUjMwWXFYOhFhQaV38PseIw2cE1d+sm6u
VxICTsqDVt9FDN0YU7G+snvSycpjMOnERyccxGguAZJhsntch1KoXyzaN7ln9QQewjyRCz+3ii16
8SbhW+T6T7lnwkWGWNn0LAAY9zzzHaQ+TuICgOxHKWOWzPO5sY0sylpBoYhKH035V7MlMarWqH3j
4s6aR83VfsWZF9txvzv8IK6s6iNzGew2E4Mgl+ZvPZ0IsnPLdTDETTle0tLN9b8WQLeebUOa/5Dv
w5FdDVZw4yx14VFrddkxYdZxtBZs6+W50Cz5rEzD5H6COAPuj9zgTKK2TTNqbjT5gonyZQ2cpCvo
NfKp8tToY2HqN/mu4kKUjy3qTqjEa9gYjpK4/exzjPMSDnjBF9z2HtoG5pOwNqD3HXs9eyFGE3io
jP4oEXHMz7xet9hnHhRZPtCZvk/2zidLVWMv6uDxUJLJEQQOX34F1UY4wq72zBYPbC37S91JJ+Hb
GLWqpl/RaB+ItHdLhcdA7aX8t5Vd1vty0e6zJh+8rrUTSz//e8G02CKVVxx69wtum9QLZjrBg+7r
71qHNykvvW+4thEviE0ZERjNuk4wVcvnGT7Z28Pl7QIMCLC6tCmP+9hyvdpMFS2RU8XtYPbXn8Kq
M9yWDpH8R2c+xENKzxd2XADSNOcPjILs+L6ZWDWsDbDOlLwFVZm/J9jZx/Bw744S6fJoZo5BKjoO
qJWYcaJrX15oSTLAH/aFMQQ9kLMQ4aJLRoyWNoGRZE7Z4FY6T+0hySJdcOV6bIi4Om0MyaoBnqe8
T2jo0x2YUPiiYqrOD+m263NBhpgAdPV3nl1p1SU7A2MXWrCNhBIxL2/WTdAbYy4COIVWK3mep/QE
5FCfmypd/Aauc+yBRqz6NcvWh0MLpuATqTjeWaakzCAmAsCx4k1MuQKD0gwFfMK//HwQwkPEjm5q
/HHiFFiNkrNv5X8JcFX7uAimut056AE2nInleCjfqdtEygQoNr3sEa6QnDtYupEzJg18nTjNTOht
FKcU2HiO1Tn40MBG/o8J1gz03PmT0UF8/S3wLRXa/TvXKnG+PHok6nR7BTP5C/3HnCsLVgT7H2OJ
UDW/fTTZdGX6lR/ElCmAEVDoJ0zohHdJRGI+BeSfywuXc8xE+tQl2wcuqYjB0mq3wz8FfiGdj3c+
DjfSV02GGXjpxNTNXiXXYtCKihgwXnpthL+owg2ezia49K8Bdk5EZaufXJ8M/WfEAtj/pVEp7fE6
g6xmlGljzDLRKoyusTTaNYTnNJtutaGDzU+NMZdf2/HxfQraBSGnLOys3a8fuq46f+v1QSa+h1hT
lFUyCTwLtQj/3E97lNwcO+NPUU3fZecm9lau5GAX6PUEgYZU8ki0m6UPGlrBo2r8GNgq0zkeP8tn
eMSK+3r98FszeRLLiPJ/b8HXUwgngKZOFyQawwwJA9maL46YCqaagMN+G7QW4+XKWzTjCb+VyAv6
4sFuSYEFpwyr1DMI/naAq12uACw24i89YMPqSUPBL1t1cIUHgeB2uxZJk/abrEY3ttpEDovDKpuE
OjQD/AK48d9PFMHQngS3d0C2icF9OhZoisN3XA5PFBiqzCE8T2xVNWUHxuGcp/r3hLKMTmOOeWI6
fK2lN2ooPD8TXhUhl4F9H4wbIjFEWdpzNOzJqWM/zK7SW9M149T2JgtYtF70x2cHhUoUDEgg1HBL
FsbxGrafx31HmFgLZBYUoX2eQRIGYqc+1wAjwGzacvKjOoLYh3kUhFw3QvPgMpJczGs6KIXfburJ
3BEyfHUGHm7j5gwDk63NgJBuOEJ0EjkI9jZoPfrU8/6xHWJoJ1E8ukXwk0pCtJzTYpVXxvW3JF0n
FkYMyTAd2jWqsyNgTH2QjFwjE992FDPGo03jGygmIFB14lzAxcFhT5OYp1JGqKy8ag1FnyGCquD7
FtuQftFjE5/l3csv2QuLXBJ18QbGyboCat3cbzi61tKpgGYTR/oP+Fd7pC84IcPbL0kiMTV4nXp5
tbIejU61FOm+Cj2zRJqtWWAPR3U+yMnPWVjjEoEWqXW+vrwruZa5zixVlJgY4AsNVBkeH4UGfImO
e1iUVba7Ei/rECr8t7RWL/k6YuAX1tFsHDZBMPqxKZBSGdybtS8PemapHYi08bkPcpKna+pL/73o
FV3q0iPZCk0TRuBo6uKCwYucuVZjKxqfJgUcHQkAqOa5uARi8I5DFTJLw22cV4+ndYChbSOEi7CA
0RYbGqXZBbzeO1QRQTJhqBThR/45hjH4ZEzArGF2ZGaa6AeJXg8YegDuMsqrW2iFjebDJSgYlxsI
cyV9aS4PjCpmNqeEepGXvbqDXyHq0HajA+o+mcusG0j/WBUMKakoUgEPXikC86oK6TEQAchceaLU
MS+35dgYzLNZ9LmNKcTdbyZd9yvCuXcogQEEQQ32EPLCZzgsI7Sy43C9UqJr6//Q0rVlxNLZTtIU
SwvMZpayvg2uErXXVp6zQ779wK/wt7yV4OL41nU2UJcPcag4VNvIzvmc27aIikmchPpX2JtszffM
R3W9DBYSA9GKPdXMmOHX26v7aBIhHOky7OHx0DrbdOMcedIORH2N1eUj7aulQCCmGK1sNhsyg5c+
ajtvhaC7R9z0vcMWBDnY6cARi0vxSIRudBPJFdXxMCYs853NKJJXxtheaWEbQsJqKQtv9AV7/Hc8
rlamgfVl+Fvg20Bjp7rH2haOXLe7Oeq4i7ahQ7xa/ppDNdJW3bY918j+TIz6qTPtKJHZQ4ET0LoO
x2DMG5w8y5A0al/xuOLUotu3aThBCn4PgErM2VjAqVyKBySnfj6QiDsZUSWIaiu6GSHKAos5+/5G
idl9w0uwUR2nXk1+kll+cJUNfO1cQgT+LUwVrnVxpw96VUv542+VBTgvmdK0C4DcNNOHWmVNoHGD
rjE76kD8X+KQ57OiuXR1krA+L9eCflPTyD9AdjFVffYjzV+8zdfb81J7zZcJqB9E9gieGwi1+g2g
6VawZxR5idbFoW9/Aoxvo07m+JGZtB33gXWxu+p4yTAydPJjEy124KVzrCRiwgu5p7HyLGsbIWVd
nH4GlzrJ1nbLH+hi2/yA/xzj9dsLRZgNSEIwPGgYSuoHZ71soSFCL/5YK48ygKsXpUfdOfcDk6ub
pjUy1DMxJ6l/VOdLKiBnXHtFXbub100CN2FtkDlk4ItQPZ2i/09e1jKVzX4RBeSw757Yg+cWkg8z
AUdDqIcZqTmtHkO08fz2b+5ItMATqH+NhWBt6X3rjjZ+sYW4Ye9F5uwT+tlMkJ3FCK6Z6K74I9Bm
fo5limg0f7MFu6ritsyGID777cfXGsFekbnddhzA4OdaeWub961SAHub4TV2lMRf49WbwLix5j3e
xERXmtLkFADnG5TLsJ5q3Axr576mKUbgalP4G7JTCc/Rvy1AescVw1ujlpiM1vEe6oV8WzGsvO/9
tJXzivgKdI7zEmtD2RWjbYL8c/klqnRSWw2NAFcTU7o45+mBrH6RWjU2b6sDp/vTwPRm1KMKYtIz
mJO7/l7+dfdvnGITfvqDyj8qRhSY/7O/YIJTFF33oQjTKSg+0fVzTbkhhr/W0/7tztfnhF5J8KDz
WpAU0Kz7iYx1yR/lGLELAbnhEm8B23bRY3k8rV4XiUiZFWaRt6ngt/UO0kVZEE0N4rUnyJqQjWus
ORPbTJktLHTI2OACopMx88gWmzmh3fxzCk55P6OGB7aYevQl8GMXC1Ac2+6vHIqwFIek6q0qrppc
3uXZaYjPuINMNk/fM2w8qK91PKanI7DRJb3Zus4mwbp1tq/Y8awJ8+W2QLuB1EesB3bo9R9790mo
jCEW5x9G4DPE2qR8O9pizbhnEnSPuEP4qFdY+7zmPF9Oyv6W49np5AcrtY18iGPjtiKA4F6OF5z/
x9CB2BtGlnBeAQZi4Pti5XCUe+TzkovsRMRYJZRF24d8WXV6SjFoeA3lmTc52ZR+FFxHdFNJftLN
W5MECRb+8Teh3uAzj33hcD4RFCTBmuBZb/w2c5pagTGJzwN2oKSRGvb+l+4+UXCwYt/HjFsEAQnC
OqCSFeBrrI4RQ1UpCfeg6AQ90BRiw0e0brwk7QGH/qjBlfffLdEp8FuerdPB9wHePpJkrXPb/aWF
VGXvOxIvtBvqUgPJTyfmNsRztogVpC2HhNXjq5yodXavg6diZDiy2xevoK7MvqD44e+qIdn3gTOx
lv92UaDRc1uTu4VUAMAvc0PDYBLqgB2E60+n5m+GQ/9xCxXSZ13pnJjKaMVDIQXEYFrePhsH1TOZ
GxMMeRXnh1SqW8vm07f0aeKkMBoiOBYd8Dy+Qp1NOwmqkd8fdO42VQArCIlePRQSzeHNxQE2Vxqe
ZhbqS0rqnCoW2hUKx9E8JFHC+v1WvGa5DHlaGN6qz6v9nrBb20ClvMmCeKQUF5vGorvZI3lUnqNN
kgH3eWMvBER3RlkTVZyXjku7YOhN6TUmBtAGgQBNzD89gqu5v2SO/T85Y0OA0vCTWvJq29ejLlM1
jw05E5zoNWCkoRo7s+lAr08YoTKGNksbNjZOgTyPt9X8bWVqDKN541mQhTAyMmbmpjyCKLLrquZu
Ll9AJlz4FkLHfxXjTF7+JxYeO8vnbFmYZ1/W9nIWt4vszlx+3LWLJDm7DzSvrqzCuXLNxeZKZ7ti
MsUbIJyDFLIu53E1tHEJQ6W6vN9+UPj3HSGv4kjo3gIE1t/fiIFa82VhvtpWitpX4DawdxdAtVs0
urI0n1NtdMEfkUmoUU/r5YQacxdz6aPKfoC6HRkO3l1ZIriBHb+Ty7U+rIcPDQ3ODxRKFUfUfHcr
CDrgGZAlQ9T6yEFEppQ89rPIhpXaiYuy3OkrfZh/Q2wMMhfl0D09EsYXqmF7W/eU5SuJ3resOV9V
f1Im/V/9ckQXm+AUHu6QDJ/x/DzPIDwox/nSdCCslFe6FcpR+KKXwe5dTcJVhi6CCGVapx4EEyIJ
TVp7aWrLAMWVzOD9qjO12ZI6Q1dVYqRR2ItI7OvXcTReAEE0aIF2XvUOLnXfTmqRb548T2p57VEH
+yOETQnRZd5j6VMLlK88ws86xfkPfP/ifEfUk67Od4zaFsKdNiCg9ZRLkMjC1k1dD1mAzfX+54Mq
k6GaSDKXrRkvovugS/nkkvJz1Mg+YWdDprJCimzkxzSu2EGPZa13jN8QVs93beQxx7of+ab9sFZb
TySvFFsGRQAdje8fXqpgBq9vbfQM0TPRpmv18yMgOx8ZPlXBnVHTG6KhG1Sn1sgwiqI9zYqVEVPi
tTTEUVD7I/FoxH/rmLan/FcuPua18pDua8t6vUk7/Ru6ufcnQCGjEYj/61Ac+hqonLLX0HzC+XHA
OaId8lcRwMnLopRHjc0qIrsz9VK2BLp/t0FPjoBagC9a+wKynO6SQ+RqvyayGafq/xlNBgf/QGWt
/UWG0ZFF83MR8j5WnCM1t6WyaUxfzD48uWPFOqLomTHbw/NU44OoqBlDCJYmCpd4qrKIMkm/qDde
h3d5i3gFA7FPs77+38zYARc9QHyM7LFGhcJUb1vmIxtdrXBPv+ElBTaevFUVNfxr8agazHG0/llr
CsEmW8iPqvrDewNKICbXq7dzvGFtmI9S7ONhxwpASVJMPIPZKSKQ3ysjCxpM2aNOZDs5INSBt6uy
YeE+Mlqo2kNCN4gbF9lJwxd6b11Q6UP+GEoaw8a+9Dwn06slF3eEjE/nhnZWd9RRmwe1PaSg+V93
rSTqx7RccFaZXU6ZsJHaldPPD2PBkt0iWyuICNXL4Ucs8vEl0ZLIxbrHlvdxLul4Ih0kxq6K1bE0
bxmyUomlJfuaqXEq7tHVeZwrHap08hsH3DcjmvfcGWEaRVJcW21zvNeD+N14m9d+i1f1p81PSU/T
towZRB7c4TwHxxAz9Zi3tgpmO287hOee3LJOwfqMo4Z5iuFPjT//2tFGhW47mO+EazSZE5wP2RRD
Pa6MNXkM3EbNHbkstTNTnWZQoLQ1hc6LpRuYhxmAB+LDS6jlZpr0GQbXBgkEcRjkpqjx3JdCvCql
UssJT/o8pQpzpfsDQRItR9qr7POJfu1Kbq63iYErjSmElTT2RHoSuk5IQy2UJcAjqcM3BIxJuiv2
SdiDDBo3z2XE7k63j0+J3H+sahwn/TqZ2f8mbyX/s8YcMzp/ubJSEiMnjCs/NBoVnTOHUnBw1dTM
7DkdT2m9t3aYI53OMcPr3GjN5uTFZVZJ21ufZlhuxcZmd9oW6qb6eSQ0XDZNQ8QKcXeFpzsOREqG
cH7uednEuD1Wga/zIMPXGoDBs3hdkeUTxiwEVKtkHhLtEdcOBjgrxlFujusCql8/USS+QNBNeAc8
C5I8yNWEPwlmcxXqz7cmOS3gTK/fjqW3GFRrb2i8lpQ1w9lGUfKTJSysXPQ9fUTGy7DjB+XU+r2B
H4rC0TbGNdkFx/RuVSQr2LWLFLdDpIKGhn+ZkA9bNwft9JqEa8UEAjefvhX5waIWImYgVbF6iqIH
VD0oX4/aazwzP/rlLt0sEj/FVnaiwV9T2wGOlFo3ISLwf23IqoT8oVwrbwz0b26FAmD62PDNoeZT
nv38vdDN2UP4/y4iMRJNxXlddZF4KcbVFUy3ly635tPSQ+Gez2Xpsc37f9vQIeJBlXT4B8sQ8XYg
Tr2PME+tzypuO2ZWjZW1SoVaYrenvBL6IslboYTL1o7CLs+2GCbF0RkRZfH5agRAGXs+7WHvC02H
86+OfZi2wFynL/yT38uNejWwmhoSW5/bTTmcYgG4m/b7yuQwVlJ4XjnRz1S0JdSvzcVPxzzKiMHT
gSHvBxFsD/fWjRxaiM8kLUU3lSxRByWGwiVRgxA7RPe8ZdiQRjjVu9W8ZIJ/cFGQ9sIQzk2UaCHf
ENMyfCQSbP5CHOlPQDlroq4JwnWW8ZnK7HKGGwQIKwOVHf+//ssZ4djWvwjgKBlm2gjGKZgFVHPr
rAGVtvkOXnqvj3Q7rnXOkosKX+uHPfixd7aHI3Jc8RkkHJFzmJ8V62WkbjZf/0MFVjUbvDaJegfe
wBZ50HLsvgTpl+5iizKVtMoxCCkxKrw/CFK34RU7IADQYXc618lZ65A2qNARJSz9Dj9gGEYGd0o1
e8d5G2N8kLQfd5aj2Q4C3LaZnvqSadoCc6dRomgK8xN+QTcZ9bbguyWZy5PzC6uVyjxrdHApedvV
hrARowg4xE6TS9TRtkI+FOefsYNhdhEY8JL8eQl9zh8VgHRgxc4ovPrXIKaXHuqBa3ua9vVnUcX5
zrnoOEEhXWsSyuzx0Vtfis+eJBlZAEmNZoAJRK7cXqQoPVRXB+8/0L8npqfeg5l+oM7T1ZbXkGrv
VblH3ffD6DnFOYMPt4rqr8b+9dcMaSE5sXj5wa3Uy84NmK+XRw5CUhCxdVDVJp/YliV6Uue9f6iG
9dgJ035VXw67BSL1GWJMYMebG64Uc4s7JROHUVeWRbDKLnd3GCCCWLCy7opQnuMFpkISdby9Gk7a
uDSAieHW4V3pBJ+w3xQ/54lgRJcV0wQ7XqgSjw9ojwnnrX2MqRapblMXcnyk2IJGExrV6DlgudFS
/Lg8IH7CI2/9Davfr/kZ3XWgSWUmpc5CVNU3faRWrS001BcQJPtBg1Tnq1ZGQtqrB8g9SvfgDeSK
2Y19bl55Rg8MmR/4wDMUqwNbxSgAXe9W4xZhIAYAouLTKDHN4bhWmXwuqglPATly9EoNjVBhYej1
qopMAnH1nH0PCM97ft03i4KH7w+LdPqWBKlzcnplbrErG43svZGu+krrlgsg18DAi9FB9xEfUrYg
48YP5TW+0LbOE9seLmnAjndYyJjFPqX35Ga/0nkXwlwrhCwyPXrFKB8hTA/E3KEMoqfvUeLXmutA
uLMtfX0/R0i1jNSkSJ5Y5zgwdJ+mwczJXZP7mJG6iwC3wthg9iJCGh5Lf5D7QAWskQSELgEmY3e9
IGZN9ZDKlStFRuOzRVkXrR6QOdmtMwhLZnPuoAQQMKupgLeKhlbRBweqg2lP3/PSt+q1+c6sSUdV
3rgN6jLY0TPDNA1FVY/3LBac2R7Mc26Or7E1Z9qWs+DBp7zhLoDsNRG+nN2dYfmPKU3VHYN91wSJ
SD+VE6S8nt9LgpkZu4/AdGa7lfJp8PwG0NhJpDVyuYZAplIdqIDTiec/yKEyxki2nXuNqq6ibvdk
Yx2eHgW+8eCaW/AgPX6tDiGJrEHUnVu+xWT5MOqO2nHdJKnBHtTxl8kPEbPOrAvW0LAd3gqfw/T+
QBE5gXuP1vdlvx1mueoyAHhaC/W8OpIUEbz6HI9kG2Pow8LvsEioSCH5A3oWSIq4hUkWPddvtGEg
Dz6j8/bfKff1MYmMAQf95gt6L3Dx/Pym6O4VQ2ue8u+wEH1W93aAOficndAIt7F2AuuXs3Lu4D9V
b90Ut/rwx1XSN0gL4YkJwOZNTpbCFxQhWTKBEpFrBKGiCbKPk6KWQ8xRksq7vHzruu2ZxCMHcX2f
U89GMGKNOgjcwQpR+quEBeUe7naDVKBw672VsaVLaqS4aXenI/NaAeMC1lVcsdcRQzBcYhN48Mak
oed/nf8z5U5X9hGApC9aaoHYgSYuvL6klB9wFnohKoMd8hamV9dRHiHDTZM9oyVS/vJEYK2XQejZ
4zeszF6lsXoZig2GNp3Au8p+LgWL4sERKyx0yXlSeDVEh6T/BqTGqxcfkJGRfUooyDHPPs8T4IPm
Nw2PjTRl1HspST5+Yb1+RcWV9/I7FjHXBA6KCxWakhvsNNrsyq9P9U+XyB9k42wAEerKEuXBzjtw
rTSyaNdxCJ0E6uzHQdB1zS20dOM3y0xpGHR3X8nKmo/2PMAFjex3E1hojOY3he4PgExXRoNr8Br/
053L0DaIvCyRfGGrE04W/IHaii/WseIFH4G2YB27Vtz3l8uEeajNFgdyhcLUgEpM5zL6RMqgD+z0
QnH6qxgp1v6WL0YmCArNj8991tOPe+mqxAaEhl3kiJhSZ5qBGxWLzRMKtjpEqWSYcGagTiwBbrfA
vBBKWqjSSaJgPsQ3b58wF1mvpzRHSOd8P6a3LvMzEoQRVWFTvFN3LOGiJNIxFnceGvTx7UQKU2qJ
ppw/SoUKi348NRRWdQcnpwAroxK3jtsROvXZLn/gnc42FXNfMqmVk/QpR+O/FRy7kRfuPAaQ7sXF
WMaMlMHqlEnqXwgwOvTsMUUb7+YwfSJWAR8y1eFvgYQznuC1QFJW6Ij6utA+4TcUQdn/z2RhJCD9
SfVwFfFa9UooF4ZnxtTrJxoTOfQSh2qwJn2QycqHaFiqXtmvRY7vXe2RFNDKHShVCtV4C9rY7EmN
VDyPEXJjiS/CwFGJnYN7nDpSxtGPNln3swgIhcNCEpndoAMhv1bYOX0y8P13xeb76Up6KqC+XN5O
NHHQRqX/965ZTzwh9lZT/BiAKV163poyKlryZXDYBdIvrIGZ+R+PTk4uAu1W8exIwqPoMIwhGneP
uTcpHWlEuhSI3ofVbhUvN1ErSrq6pQXZU9l/Gncqaej62PVJl2PNplDOFw2i8OjtADiP5Nx1cHWz
6ZsuaFhi3nG4D7hUBbTU1dxiwuCf6+351oT02Mz0hlGBMp9/A6kXLimV2JhdGrP3Nyiy64FwYpHc
Q7flpWy6hK8cDVOaN0FbTW/gE0uIIltyotBQt3QEqm5aqZvbSQ6+9yjqEEwAsko+S1ZeplwlstF+
vYoR34ZZBQnwXhYuIpEH0tPRdTZyIXZ4W9iJkugBQAkMI+On8IZKI+vL4V5ztcNb9xcAvkDx/4DK
V2UDsIAgHU7qAro/T0hur8bDCCSuoZT+nzKYybKeBceIutSYif/YVGxK8EWhsx6hV1EujkdGtQci
Z4xP+TMUL1xs1Aknz4AF2dKwrmL41lvQFoYKLRrkBWq5sIk3w6ndmQMXY1gPBPn5GgkLNRztZA1g
eW3m3tJ7twAbeK4YPt1jIAQeIMc4ClGUw/oBTuHCOQ+g3TdIIKNSPssNxEyUv1M0oDh3eDuwtxM3
z/9du7QumySdFTgozYh6b2Mv6+zlbRTZG+1yWZH/3idQxqJCiFx29J9b9U4qRFxc/3i3NtLUXwZG
PRKAFsaI1wqmToOg8yKTmIJxRSt3m5NlLqaqp8+iHORcueWeYMP3C+WUUgau17zp7DYUBMptPTGd
nlKW6Lk1YrRynooh0EtKwfK7NdI0C4wh3JZ+RD86iYpb9UjKOoirmVbIYpT4KQJDBEMx6WUgI3u6
4efSGkxTrbouHir1gc2Qh1ZMwykG7b9XFSL01/qWAD5JHxtd703dyMG5o8T4Tfywwi/cONZeOduc
uYedlHvgBWct5T6xdfELRBIr74KOfPYoZiR5s+/McI56dXbIfRddT1SzurUQ5ISCRWpqZDj6oWLs
UZBajbnK+J5ti3BCla8yTRm1Xiyd3LH33G5y/TREHrL0GzjEYq3kL6xvM0oSMlEdXP3lLsAjfyKz
p2uqlA4VvDmzcnLQWN2wZIGlYam1/eC0pjD+8MMdBJYnKDau3yJw65u+MJJmrAJfSeohs6jQA8KV
PkPfkPUZVVy3as3qjsdTp17i/mHp1829llkfe2N13UjEwVFgv9SXvWc60yMZPbnkJ7Mea5h4hlAU
D8o+XcuxSzgL9Jjt9BDvMjrlRnOQORJkK0AarIEQpszhv1icQbI6B1rTDSsWR0It4T4amFLFgbED
qVCTaEbSSXwckf1jtiSZEsx3xu6EuOSI8X65C7ZVnFAQ3mhFTHLaAMQwNjpHlg/S1YYdHwXN3RIA
fBIqccjOIXAoejW/2L562V2KXc3l4HmupW1JQgIv107QGhZvKwVU065FCi9Csk6kiWGkQTB28xF9
MGCNQ+yCNtCbxgDnUg5Oa379ktO/17LWgFwYtJ+eLf34p9b/cA5DMnrilqMCFhFOU/MYsbMopgbd
yrXvs4aZ/rnTR+Ej7N9giiwFtAESZ5GojRgXu09Ts7e9oJKlrPWQv2bAZ4rJaeDvLM2fEJ4XCWY2
RQkh85RHaHZuEysxU3ohKJeFbz1/K0Z7OgVNu41RQ2qBkT085fHV4/AbctKpe3ot5j5BNEEawo3Y
DFXtUcxbTm7gXr69maL8vLh4Hnfq1ZyE8on0IezZmOTSnlYzhvWfO6JdgJvJcs/M8YAYV/Pd1SUn
i4JKEpVcQRirGh3P3yZDnGszO26Z9sx8i1oyisvml4wHjI756JAD7k6L2IxfufB0JtC6wOLLKxiX
h4GD/pDI5S58QcdfecnCA/+QEjJEWQ4Ji+miWTRnB/usZi8Cr9cHLYMzNTcxdQGq7zTy4dSVwtFv
/QtHAb+zmGnPFUL1f5pNYRiIGXPCvCGRaSU2mdE/ecLppi4YIV9VY5KRpRM0oP5c+jNZ8qgt/U1K
K1rslBt+oOb1yTkB+ebqOBBqDNdyQqUr5LulmRs0p9kee4Bh7PW3URtMW+9XC4Sj5SAG68z1VJMg
DYjAwFu8ibneILUWYiAd+WQBbxrntUB4k8c9lpZsvjqyW7Dy7YOxuj6OXStX38N3GEHVfnSVPnxw
QVAlhsYYxTcNevC/J9LSd0NNl8/FMx5oEKJBW2jQDg54vMU+1w8sQ+IFpAaAFLPkuPsiMp0/ci1v
kBkrcMGoyyIDVvNqmtzVdcMS+xllnT6LQJ1HKXeGqjsQGC+IxR+BkPCUkqkcf435xSKcNb4Ww1pu
T3xM8let7wvK7YUHKabvI4wCqrBUrrAqBZdIaK9G5tu+NvAJklCrAF18YaIwY4ODcikfVqIrnNcT
1CAdjcn9efhGWXgw5Jnc4jbhApPXrH3TXHIbrytpJN/z2cuQJFL8Azu6AZclHYe/7APiNc/Zj9oE
cybV0pg9Izot5+p936JYDQXeJ6KLIDdnuAwEMLo9QeeyAjHholY4qwn8MBAtzPz8zn4MAiP9NOXU
xYXr+vLkrx/dHKuvmhwEYoQRSCVmGeaPRJ+j7E4D829pvUifMMQ9ahSOpIybASBje2RiSDoCmlm+
LlaOFSJ70msfvZxRlsmcrrwoDte3i3qiQyz032kcYO5sHchs8M7N/FGdNugX73f5gCp7gyQSrFaE
/gIZPrhVkehVqr//drzYwBPzLqIWhVsgEvJGNIvGV/IFMYbWhtU5eg80hS7V0kG3GjWrkuHBTeht
j0mm3i5pgVaN25DvJMw4agDTIYl1FFW8279oYANINzZF4f2Hwk6iSwt64Cz+91+VhDPXYzZQzdsV
VQlxK7nipEXnTvkPgWF/DBb9gYPZMd2CbodhhgNtohwL9EY43zQW++sD3dp4u85kCFQzZeqgn3gC
Js1XB1t9fNCiSH9GKV8/0h0s1P08TpxD5GyGheKgoGKiuX/o+c7lN8EQ4z1MWKTZ/pdARAfDeZjA
THf4uYJDBTNVr1QVzfImdSfVBdoK7jbsG7d1jtjW9GK8/wH7OYlr0huNpJKLfGxFmEkQumPXGtbZ
J8XLomMVvTZO/ow3AZyBMOKk9jhkL2GqP0IMrjLl1L6I/q8qP79eh1IK1hf9Av3UX1MITu74n07C
a0uFlYWU1ZUH8DXZ4YoSSwSRPkxwpm0Wp5RBheWDpgn/GAYr54MPVioSITBBpPY9thnU9WnIV+p9
4CGEyNMPeaUPQzRm6lWRmRhN5go9/AiyFY0U3mfqreY+jm7EGXzufQoVMR+Nhb6kjQ1PuaNvTk8c
774DWbmmsWsaCI/aqYOGH6FOW+fBbsKcaKLyno2XTGYQV2PSOhW6MYB90RPp3BhEJvTYENBiwQ+4
YLtLeUj+KUO+EP4TYDTRg896AZ9ek1Koa8uXxJry1JEM4m6VRZfKZRLJ0qnGyvrpu+StPiykw7NY
wuNdzW7USPMStKPjfeWeIn5EhdyvAS5rhULUwB7rWhMlsMUmCD4kpc6kwdKJ/7UvMwMsLOq4Yu0T
pYi93XjxY/lyTjPqpyk3IW5Xop9gHP2BWuhpXOMnzMyBs1MOsn3DsgYkuPQuTUDjDIUMtI8+4Xd5
kDnKq4lYFRh5hW774FlpMoDue9BqCFCkgmpN0giJeoES69M8+2P2/5bW8vbZ1YQ796yXe6gqLv8f
ySjLIFoHSRsgpXu/bI+F0mwb6m8PAbm7yv/P26/AK9+ICSH9DfZEGWSSeMB2xCcNTUfUZ25Cym+y
L8Kqn67L1GjDrYIgFlDDaJc47GeHZcnIyY/+Lb+uh3++L7c3KNyq9ul16ypPrJ8TCQjGVPhhNeOr
Fa6QEl6IYJgNzufAI+BtwNCHo6d1MAGqSgJHMbyVA59TYgf7+EYDfWXWxAuAFx3ASOQJnt3zE5vl
rsGZTo2r8WGLQ+jeUa9BmAyrGlkl9Qi3DFElu43fJtYDG0dvs8RBcc/VvekMg3ywl1KvDkgBV9Ix
SNZ+GMvYVtadW3swZZSEE5Z0tBN6+HTw9f5Imrua1CEDRiB9PkHPDumCp0fXpcCMmQHgmk0nx1Lf
A23oW+X8H3qniSPdN2Nhel4e2Xv61DW9abEdX3FZzQIe+fFevyQ6jnJcU4BHws9xgDDYxOA9p4hq
Pec7nP4cCVFl15LZJdUy0SZpTiFVlYTkPqi7ODsOmZPQlSZekVriRAZV0Ry3oh6+WHKGUXgVUU26
hUCywS7IOY3qhZPbinS2osb1op1d+UyYzDkiRkL/pbwOqOvPCCFG56L+B5zeLmG8t6brlroFsDSJ
JSU0+QGJ4GK7s8n4RpsTvKBm/MWaawfP/w5E8yR7gco4AzkmUv0a1CyEqANVFhsRSSmnc2RcYPn1
wEKUlwB0OWw4PF+/2cVJi3r9aVdvTuEslWDsiNhodu7lxHw/TWDBzMmUddN0J7pUdcuD38kJwEqD
SLOXxxQA/rWO/MyixAfmwasZrxl6gi1OHNPGQCjNxy86L6s6Vqnm2BPDyB8lZ7J97/kzm1/O68jU
tR6BqyOJQvQPtn1eS1ygixpD4kPhm4uRG+3CNWOJMK5E5qLnWk/cXJ/U1v+B/a/6cnZzFNzptE9k
pQMm5dMBz9kw76sgq8Ih12f56C09MJaBrxS+PWOmIgb8VoiPVMljDSQBpYdXok6VxZzAMbeL1ZlF
MVtFLLd9RHrViehI32ReloH40N/DWejXg30QEhkn+RrjVW3Udz1cOouDeVQjPlmIEICv9uq7Gtsi
4gMmPI/v3oXTS8Sk9RlkzLGs4x7algkQo+Uf9pdlsLhxcWA/QZ/W4zPQeNUY1aiOBW7EHaUrabXs
KYvsavnwOwPMONwisAj47AHclQaBgK+hMrPa9IVAP5SpYnh4SLmMnZLfBbG7DLN4ePDrUvIaZegq
UZv+1FOsRt49HCWHSbCc04QuDzygtU1+SY3AaBFmKz6RBJvlSP/eJh54zZqy2tA0UTm/96sv2Wkn
RuimxNJrtO19UcEPgpiW4rDCZ5bB3IPpiCVyyGhDjZhQDj5iWncTHoKcuirMdhlOy83Vkgg8V7Ba
rxyWFUMqB6/e2vregqdaZHtPVSehST5aBm/h7PdPUbFyjhLYadtBNZ8GXVU1iPmxFxsZdDfiSvr1
9I3/NUm0b4jgANfwOuyMfFGRSFapaq2rDlypZqNAGxbUvMFOeErfvGD+p09HyumDEbDvxy8dgdUS
RN8QKPjz9fiw+YTSXAzkCU6ZjSiIZ/oLT+CzYvCC1hPlO2QeoaqoG+PJg0qFonjerxEqtIhoZtWb
eUXFU20B21ZxI1A9RQxSLZyasooOK2V6EvbMjpwR7U09L5atO/mZQrQxol08xxKxaM9xRGgv3bNb
QAsnRJU9QIxoI+iP6iPQLDGfCrkDMQ7vD4t64aNdLCgtbHAZeRdeGMFj1Sgzl2HA09fvjJn6gxNb
rT+VF5P2bSgHRQSrm/9hqhrpvWDbVI9LKs8/sr9rJ+u8T8l+KeHnIHNPDlH/BRKwEuAwfYCX9uev
hXYYfqLv0zXWDi9EgREdqfnrwGXkez3iWS9mQRp0EvB8euycUfZtwxjEbrCxFW8fkcipUnafvwyl
bdRWz55i8O8wLa36E++GKy1yoiCzJH4B+m38yP4IbPoPryhmQ2gPRmbgYkCLVrBwP9XFB8CWlA+B
8Tq5LtguuhTev3hm6krVqmyQgW+9gAljd+th3XTBoAr0JguLvVSlmyicyijkBbWQ+B14MdkxdvoO
C4j964YefhE7ySZQY7DZCc/pkO3dtaSuplW08PSBY3JL9ICcvHf17Bsavuil7z30cgMowFQENLzb
LTeLfKWyyibc4P5dZ4sYWqe7eJYdYFjWOXjLVtYGWRsH+sfEFQH7pZQOA+VCKo3+gEPxyxjCyNi0
DL9iM+fpCo0pHaHDbU60XlAQjOOOZRg+fvByQ/TgXfMpEBruVhSw5zV07DpkSqUwH1GAu2gZCyug
dWpZY2CKh3J0P+Sy0cs3EZLXZT3lr1kJmW702fANoooenq84pAmBlJ/01cdMrAiUWtioFpRQr5Mm
Th06iQ5gt7fKbgoR467X9ux6izGTuNOTwXxn+5pTBFfHXXw95kQr8F5aQLLWaS+llgJFjL4YBXAj
nKF6vyqHGcNdaKuFMrFhnvtjSFZpeaJTwY//KXPJyvWb96XYJODhhBN/VaXuQZPpnlKtq+kXk/5q
+qHLZF4OPkNMu1tIsmwztjGBmd+MvvUbtCEvl/zO1wF1a54sNEduVER+SHpngtsfpd82AGECwTVT
OKJAvECvC1GIlYCowLa6jib432s7Rx77kKgoyhsGRCLYFvgnwB8hf1Zn8l6ISYAMJ59i4Mtdto5f
ewGxN2VZI9okUfXIC7and2dm4UoJZw3p69QCPEU0OFxOKhjqOK5vonLSnClIsBTvGPaUfElHCHZC
bmi7MJCjLMn1A/X7moP2sXD4m2X/eNz8mcadzOL6OoK+uUGe2kNfZDzhfXJEAgvNMpgfW53HeXZZ
4jvJHsZmsEzpHZ4YSYqqBdRNlelRZdk8F4t1ExDLvI2yRNJSfprB+PSetIbrTYPTOFNbgR55VJYy
5tv07KOLQ2nu6Ofu13o6PmJ+A2sEfY6AeJWTuWYxlREk8YGrE3uzCEzHeyG1/iyQ4jzK7eXdyibB
WLMKdYyNNbv63SzXOyK4YlXipEQVVnu3DEFUKBtkSWQunxiOjDcWeU66mw11wTOPvybIG/OOEHzI
1HD9rt1I6rsFP/ujpQ50INNeqbk5iV+TrOPEBEPAu3NxZ/RTITAeQvoSAsW6HLXmrsTbkw2FLeSH
Tl2gFHxQv8xdTVAorGnzXE3sZJ2kS2Y8d6fWAnYUXNSuxVowwUybeJhVGAKTET9094SALOif3CKm
ztQH6MKra8VDMsjUM13y5eibL+WQ4GA8F9dJx6ATyd7yrGVkiARiBIffEgCtVEi7W4DzQvhhdYVf
XzVVluRv50Ot0VAajUw3QrkYTIdrSWrZbf3OABxzJPCH3AG582gVFPUGlaNsE/2+0Q/cHXZ1T+eN
y+sfGzzPSv3WOFx80FwKDLV7bsa9wONILpnJbVBL9Ea2H3U0eKfjYPBc/7QWGbJUfTob3mqvKyVF
QQW9j8E8rpOWO14hHCD7aPGmQcmrQAc/U3s8uFhDgKXFw8O4SlPR0T0F0N5beFoxQdHSod39SFL0
4Vitj2Xb4S6BU+t39wHrIT1rEibVyzwNQ8Zr2LWAmosel6b1I4A1vLX0N9ksRqIjiOwjRhnQryW+
y8mP1Lcnlq5aDqXWUYPU6uD1VlZMXCVJ2ZzknQSIJIqyg4V1+h5fX1zU2ha2UAggaIG5z7aIAEG0
96u/WmPdb7qP2TGbClUkYV+tEpQSAxgDjaBq1f4jis6wLa7qsT1GgdWcBW/b9bENvq2Ud+C/06uh
vllu43T8MjYHk13dQJl5iICxLbiUxa4/NbSqgg5KdEahoO1IAeAme03KX/+qU3VsvBYz9Mkjiyc5
LKbzPoMi1w1JnFFi97GeBV2ifVnx6LPwQCrfqEzSsgA2mv1nfjjPdCJVBp/2Sg9+icCp10eYtg9/
xOmQVcIfl9sF4o2RKZIoea6CE5oOXjSj3F0ui08XLCRXxUiUOPZ4tL9vMbDj1wMulu420gRNiWyu
73rB+TpRbyXpzSA6mgBBMJKVzBPYZlYd8dHLXDrnn6YJSLHCXBvwogyyeCQYHlsk02R791BxZlCR
pFw6gcQZNxgviw6Ne3LATbYU0dy+QegAiPMD2/TM0Scth8Zg9WJtxytYV6BkXLjIGJNZ9juyM17D
K7gyE1/wQsgeIKjJ6FjDBwrnaGCYQAU8nkWfaEuhi7UfzjCqy+ANLo5qg5jvmMB454SlLsmxEB2c
UKvVwiBOh57Nh1M/NfICOhkQqWKj6aNGDEvvHtcVqXu8KxONRKqwdyvgqJ68YEIuv08sCSMt+IzX
69aDAK4Uu5RuNiHgAO0neVHk5YOb3gBtQqxGbup0taoBfyT1av1Oj4rdk+bOwqI0wenEyB421A3/
6YWfmi+ayFH2d05SYqVn1I4LeDwYZIoXxKBXDwob8FvuSz0FKRoLTJZrT0R6Rt0MOB9TbFb+y/lu
egTjo/vOWvARg/V5z5mP/UNRsOT4+zWJCnMoUCNo9/Yoq/Kh9O+cAnxo5q0qfyH/+gAi3zX2NEk/
UknOlqtgty89R8UVLN6wdvhoH7Oan+I7Dw6US9jcpclufoYCoNDGZi+rrqSxNEMLz4yiffAlV26n
sntlsKOcsGWyT6Fblfr/VmcvzuUNIeoG4AaFc69SnofpnNrUUoou7Ge9NyS3a3Q4bpeoZZW4AON+
RWfBrE29oeRpWVJRZl3b4oHykqRUKjMYKIKTueYj8jg/gh46phnh3uDTG+P+VY8eovB7nmSPhKFZ
wlTdEWStH/WEirUadOuHeNNXr2byrk1GjO6AAYzN265Dv4S+UpNxd8bNVgH+K1DlJE74RvT3ukNW
KIc6TlvX6qCG4BpKI2AJsrjo4kf3fetzhjJizgBI+xYGkXl2MyCYBaRv8IunOoK/wYa6atRNFKBA
LPbBC6JVs8kocVfDZ/+6X6CkvVDukgUuwVQqyodCupql/fI/2ZWbMS6ebivPv1KrH5vQPMbl2rRn
BPpK09iLKAc2/4igoUnRU5QXcm83tSUIWP71IKJTFGABe8OJVr2XAv6oh3ySVETk2KAYn/QqzgIK
f8fpXkC5Rq+qv6KO4oJpwMLrcN+IKZ38ZsKAEKQDRUkBi9SbT9ujuW+BT7NUt5Az3GAWSgyssL+I
I6E/PVj3euGmrX8seigkaE67U2B6Rq+isDoSIlAio2wUAoAd0yVagbxtvVsET3uyQB0GoQ7n+d+j
ftvdpwAmhqTMxI6ZTLN2IYDiiljQsJcidA6U/MKw5QNahmDz0mhHQkIgbQWMf6zXCU6u16dxLHVA
jk4OAujsYTrU8o4thWBFKMTkMfxcOQkGkZrrkJxF8PtV0I6DFcdWenQPFPeFHHHhn6jzYZVGV8MP
zf9oCeFKVC4d453co9rXYhGI2jWLiFENHf2r8VpUT1IWBFY4ErC7chLXoRA3j1cJPUQ9QN/bBw4A
nChFfvmkjKXM7pZao/Mx+UuPPPPNPYs2P6AUKXhdNvtBuWp2q3/j3lUqBZ0Ko6Ye0bvFR9t0+YyQ
1XMp7agF8mM4U7YBdms0LgnBa7tjcc4yOUfWVepMOICtaf19np7M7Y79yv/UPc8eshBZY3WgFUp+
bjUxMpr0TkZI27lfl3EP+xajZ2SYmHy4iM/7v1oSj7lt7n2VvdUMf0rX81q68ilJjkY037ICGhkd
Tdb/f9McBBGJl6zEMRN1Nv4afo1Jobt0ljiKjOJnD/AlmFlYiGIWdiSt+VX1nukGqF+aZnw3aDoV
KKnBS1rwz9ty+L0KFHxRvfhnXfevtDMqAjYdDt++1ePuU6bE0KtWj1Ny5XWUGZu8H28Q3AYKXxT1
RA4Pu0hi5mEHhBBagKdUqAw2Sep74G3cqxk1J48f3j2konSYnaDKk1lTujLPeEXLycWxPWy3ILlo
/uzOwLgKAfPQ3ZeJnE9HT/P03IdWW52xPmgsn4usm4nYeiLIcV4ejbSPguBht17uBQAI2/+ks0aR
y3giyWbzIf0Xy5zW4XiAz8QqCO8ho8swOBPDgHMa+OuqoCZaI9TPR7xDkFh9zcOkUAGpctDUO4qx
I6qE7Fd3NoM1we9drcvt80/u47bzxf27DiwKWljgi35DsOZ9gJb3EXjvMkjZAsDMz0rmG2lkIDot
q4rnDWX5AsF2r5eQQErq4ZQnyliKAoduEsoMJSBIFRF2A6BJC6hAgM+hHkoxMFqvKuozQl05EIGx
mGXKaBFQDEP8npApvRV0Amy6cTY4RweqnPhYG9kW1zLA1fqS8/fF1ZJpZ3DX2EnooouZbvbP90iR
oEf7RZFycJ5xowuZ0V0En3WMGD6d0RPi6CazBMXti7t/4DNWajuR6OZvNELdeyGWumPhjgGnNyQf
Z0jchPCQsLl0eSglChvSYwj1R1LV+ewaV5ef1oJuBRczO9r/haC5mfEV0l0/zrWsScrod8CsF2bU
YdBppL/JfvzoWY6P8eXjT4DpWX+oTsBSDyOGO4zps+YjG1SzWodxigdLnz9HyUlsxhRyXk5oE9ly
Dkj111Fnfcp2z7hAgBr8q3pknBJsJg2juv7UM9V6eelWOOZI7iWWefAroDGp6pN2h3JeINYaJkjY
V6zcEwrIbp48MI2PSekCVJFXPtzAURHeHArDbZI1V+VI3TajEIKF0n4SbJ1p+m3pgFUuYHmhXohK
ZgfGhr0SnGWyAwx2H2wMNTHm4zDz1LiRoKf4zKUvWeBBOzdaigX/+xBlSk6uZt5rJbn+xjWJpMIn
ziy9WXpq3a1/z0AL5/yWEvU4a4/ixBC/C5KLJTOZNoFQZx///gIFK6ivpCHIGhXnj2Jg7rzVa25z
o5s4kUZsIUa4V3bsh2qBGjl4SHH4z4P4Nc2XsqT+zvF2ylZcMB/lWKGfH/zLI8u9RWE8Vr7HoZmy
GRgPCnCjFI5Bjvv0RHMqnr/910nS0BNo/nyMjZm76EZzHlv7g2wyub0izup5OTAdn0T/QmqqG6CO
50RmUBymYRKyB6auBQ26qliDnFL/l+1FXo112EwI5XTSfl3dHbvCytqTstTkOL2ITPrPxdMQzQ0H
7gs2aEBHYDyLABDylFWaa7yv7rBSznQuzitelelUPqlxmNLE8IMX/O3QKOIOhoe9reUz5olTf5M+
N6D5sF1RwwPttnzEAmNNG/PeHrp/DhWXiA4Zfqrjyuu7wHgMIcJ15vD8FCcg9neFVG0Pq8Dk7uOf
JaoaZzbk3fffk6zxmzddgEeUcNzLGcKQ7T5RjkIwMcedJrtLrHyLJqUqAiF/HI6T3EWTC/i78+qg
s2MzKyoFiJ/ZvIV+WioGp9T3kR4MLFO1/4UQzw3BylmGHqy1JFB99lxYg+3vAaKNC/7sYbm0y+NL
Wf/A19hQz6c9xqXdgpJeqEfrv17EcEOKdoJVqQb4StZoSyuBUBWs/5zr7NgJLnHAB7ze9CFV6/PO
MFyW/1gO7s2EldNjXxePCZWNaDnpOnwAmCeu8rDSraUMpnriD9lPHgbRIgVIAR350cXHM09cVmjn
s8tUoHDNrdD2rLBwn6ZCp0jTqaRzhx24cmQh7odxf++NGzR79JrHvvHKVeG7mf+owVvB5DtkYUXJ
IhC5juA+Qn8G45IWvx6zEQrzpr5ZyL09/TxB4H2R7RhfDoddk1YLfwvYpJFWOnqLU2JRXWCoAMM3
eAav0jb3w/J/0DM8rTfFe3GsyKNfilC9UcS5sgYw1BZJn9Z03k1HfhGQJybUZrrRT3dDRdeeOYwA
hOnv3CQqjtsvQiLpdvBzNqDi4s5ekZYDivvVOg7HRUj5QaM7IbI+nd3R4CsM3Wxn5thoK5Y7Vs7I
feSazU8cKs1fdHQQy1YPq3ItvYiQKwOzRn0wrb4o5I0xUsmbP2s5Fkz6L93yi10nMyzsxlO0Hh3v
REnPeuDzKyGxU0oyOuPQQ/E81rV3wKWEGorl3H+oGiEChFbtNvlPWxAUlqkhXY5Yv8QgmWyFnOMb
+v00lpYLhnd22U5fyMjtTuq086J9E7593lMFZRcYMfjZ9rw5V3ECzqpD5de3g+SAiwTZRlELqwr7
vU0bu8pdjlgKOEBoVrYCmhVxW+C2pmoODsVt9WAZttUm95D1nNVSHtKRplrwyNvb8OeguhK/9XYg
8Cd+tQGc96tMppwaSdgoofNGoTr4OiLJJgkafebohg1SVXFCKl7x+0uysueG+PDBWRk0tsLBXtZ1
WubUBnEpzHP9oN/FFvQNBPRmMnKWRCEMguKZPjX/RR7hi6Xg4dgiEs7jJ7GQtMwkwkpQlInJ3TrG
3ZijZ/A0qTRAvvr7gMR7RvBJQLJCcwSyuWWySDPELd48kUy/RQDxHfk+ncBJtfZ0nytT/AmpLr4e
6rnupXvlhYGJ4PTiy72/bjG7NspZuUhuQRFQbuSyCWu4ODvSMXWETa6fBLGLhSN+eJ0RrCpgT2Ej
N7CxeuK++iSBr/FVx5VmiJvv8kTqseeEoWhasS0F+pK4pf8V/5RYb9UVkWcvo5wKIsmrY7M7RgZE
swcVdycLMnRKSHHF3hYUnmQNnzOxj4dWygraSEOmqBZDlEq+y+Qb8MunGivPJMc3w61Y0X2uyYSv
iHBlTK408e5B16gva7d9mN+SQ+lfpsbBY76s3LfG0hUT+aR2/RANf/+7pmDhycMKVwO+t08ccZ+2
K11Oy4W9wylJ+Vw+wfJRfx1IiU5FWIewN6cc6C+U80lkYgpSunlwryoCT7FBN2a6HYwvffc9U88c
Z0HFkbQyVp6DSJosUeXqB/P6Grp+RYok3WOy1MW/VCf4ZKphAVcSGHjttLRZTjA5ghIxDmmspqnf
ScbSpKjo4L8mNtNHBULvhnaROwf1WVq55XO87PdHzD7ALyNGkJB+2zQVn0oy6k57hPAHwytSZ8EZ
dp7vHdcEqTkUMdBmV9L/OwtTsX9HAk+1R9vXvZt5uoe2BXJ1a1G/TUl/IjOi0CcqJOXPWqfpLgwJ
IHsN3Jde8nZM8pzsHyAKhwZw/qkvt1/6prkOxfCqxyhdHijoRc/5qJd9ORAD+rPCbDK6EV3aPdMk
7sPdoqFI/eZifYXlV3inVXAVBpiDomJYBhOlYcJfUfhIrPpSHMi7lBBlb3pr4/wqbfHVmNzS7bXF
jWgxjqHyZnZFGYYrEVNltlU9q1JLwv6RmO/MKEPul6uKxMKUYVy8GkqwN9iGcvQh9jhfR/smOQxW
bXoemOjN1fu0y+XybrBPYzBag62PoGdrvo0IymFXMJm10gXSw7coAzBPcNdJXrQCPg0T96BesWNJ
7LYfyId99K4sysICOz81NyDazBG1D/YgJKC9mdcn28UJJMKjDHd56LhWl9cvVaOGT50DC5wk65qs
W4XB5fctyqapLmd9RQ02rdcXFX2URUPNuee6XbQW/uZU1Kx7nW8UTrdhN5Z6+YADhCJyfZ3/37od
A4Dzb0KPCqXqLmuMk6vVFBYRGTHuq/Vtia9ycn9sCASHDHNdqfJoh5C5mxuv+SV8p8fKT4kr6eDC
FLBqj1s/SjIH8xYBnMIcxvbza+B1su8QYmGZ1BtPdvouwbu86j/5y+WsP67/Ih3SHXbbUb2EP2bj
MNbFwlPmKip7SyB7B9BK1rEmWhoXCcdnffjAoFdK+60YTIfGxaA1XjCUihAnXFTXg9mbv4y6rsQi
7OLoo0Ziy5cdBLV27S2Y8KoEb2d/o6W4uB87ObXe0+rQboi/6Hz7Rs2MmrvD+1v+diIfqufFeMrI
1czaFKHMAbHJPHt6SvEj4oGEtkcdYSq1P4USV5Ac6UFGCZsUOz/iWcQDviwnzlpt3naU4E4rr3c9
JK0mUe++M6tLvzH9TG0JROi6lse7Be6jDqa0O8czDiNPtOyee9y8kfqkVx/XSpNo793sq+gL0Efk
Jvt8KpP39NYLhHtSMsunJsxSjtGv8DdPThvGQS5WSIo1I4HuJ4QXUFWR8UkqBWPfcui/GUdeDJJc
DvRYK9s+OVeXj9kK+kSFOsKir2H4rZzBQirIx45oUE5MyTnKoykfCgla0bLx0/2jKEi/GXTGZYxi
zUaDyzJtCVHm3GnpQHRBOqCDl0DblCFqr+ngPQLADL+Wbfc1HKIfLUSuklnII3Q6WLm3ZVKwbw0y
/BPDyeVQEhEnvKhc1It/ts9SIVAtigfB4b7tgJzZNIIwBm9qTVxb7eoVdwO61ORz1vePPPJGoZeM
qnEg+6gVXlq6GSAQ/V26zDr7TWFMFLzv06kolt+5jfAazGrNcbM1s0+Olvq17iYEw2dwWA4RrRVR
V0a75sfkUXFSHMtsLLjDL3g0v03S2MkpcO1gIAiSBTLf1n+uPAiL6NX8q5XD7bVLVWi9Pdcoftb/
liyfzBgcavxHiLaKp3IomwVfhuz3VbWX0p3lAG/Of5v6J5RKFTipxQBiBdbnNxyDht+Dfn1yr4CY
60KuvV3Zn70d3jgfL8Uvi0pH0pQmAMsQwQo7z+yYeJAwGW5jPQSxR0G+X2TB0tUlBWQOzG/SEIyM
HnNlcIwvsG9QulMl3BgFaoZGxkA3PZjsqZrEqLCapzH/8T0wJbl3Tv5ctiB+AGb6qwDR+TLgBqCk
gFGAbtUDBmS5JdTZ+bZyWV1aoRq3SFz+VjuOh29wBTWJCwwSWORPibrYkNoiQaNamGT1O3W/EkpR
J3CQ+AK+xtYfqyJYgNW85C9BbALvZ+uBveH2wLAhojdNXoAeqNgL2thgwgxeJk64gIvnDHWrT2QI
VX5gNHfhpbGoXHD/ErDygfAeL2qeaaQhXuts7Adug7XgRMo0QRseibXH3CumOOv19D8XchvliJOL
w6iKsl1M9FIZcNvrmG9BHd3sCJ7t6O1rrhL0sTqL4JMo13v7K6Rw9h1nhSUEjKjHJSIUkOEY2AKZ
BobD+y9d0rx3YPB3aRSvUrSfmcS3+mmAOdsBwydYifEiqJVCazAE4SBRkLpEk6Smof+cgky/zEF5
EisS/tBJcXxHxhpgIFU6/Kl5iffHTE7piJCRj7pN05dYFFrtwmfMUm8LzuHQuovuOOSQCpY1iEF0
XBPADo8mk60X3EHFclDmS1xG+42Jv+LH2EhYStgn+hsrbdKgk/2Czla8cDmGsTcsLJm6gO6Y8xnv
8meGKQI+NMe+AdIkmOev3cgb4ieGE4VDHcOHZmCI9TqMWCLJkARXLzOcsG4jRmKCiJnxUUAwHqml
G4wW4ib2ABVZigNZ0SZz7ffikwwHPoSWs4JtnPiPQpAsk3Q5Uh5IGv0MoAbMJYYHzCHgIQ0UAVWX
cYfiOfwwFYy9mxuhn3HjDl2PgSnZITCOh3YZR9fb1Jc9egmy52xFByb685Im8vYgzm9ydqsD1DDr
qMgQ4iZrGo7EdPmcBnFlYGaL95eaKflrxE65NA9xtoykVxTD5cHez9XX3PGXkY3evHMVhl+JwUfE
5b34aX3PaweHVxOsriH9ou/SRQ6/UVpHPz92aqy72JdEwdk8F1cs7KPlmjINdEgxk9rhobZ1UWO0
gXGQqDbyo6vksXwlFpKD1i/V36b02+O67YrWWFv8G/Rebkt6bC3g6Pm82BVyjecg7kCZi9xLgTEs
yWHQ0HfxKg0MG9wWRERe2S2yF3vFf3KD7N+IIix1RWRF2v8tIXOW8LkcBkeYLZBThKiSlBnGp6sP
LX8p4rzFo0Cx8+IDdOPMtYckXhOxwHEpS5mv/+f9Ht6Plw5kbPVGDvTbpF/DBbb8h/FmI1lGNJK8
lDrraefHCp/tPlcLNLBnVusI0pZA/UJhgpbsuduE2Bgd6Of3k5phjmnUKKdqhFTGmQxt5JGnJJeE
QvfjmRvjs31jqciah0fYcti9+PxxRh0mUmTE9mJPFM3Tn2MTXoItR8NzKcM8jdf3pRiXqsng83EU
JPMcgm7pswFaWU1Zwt6CaaCRxkG09gJ+39J5mzS+W9np7b3c50Molr9ZVa4Lzl/k7i041eIl1mcZ
/zeeAhF9qwVQJCsOWAcvqP0yQ2qkEqTYMC9Yk394GdxlZ2NH9rRv/IFLayRoN7fOguQs/jCMBHuB
eeLp9k8Wwy7ZwFeClc8Q3sjUlF84s7l/JWgFQhpK3erJUiqAiJoQz36rCp7OcXmR9/axNrpm+VnZ
q8Ybs1ycRriOnKVlF00McS/Rv8xBgyM+ro6OAgsvbe77MkkGchTGp7+lQ4rF20SZIzBo09R/kSDw
Xo6cK81XNRMeT7AS+ctoLIsYbMpjEpLpwY87mO+ll+E076sfP4Ix1gpy26PrEbXG+PnZ4sO3G7b3
WpO8Xw8MDTbUO3aVSVsKQwWX0/JIlT/FXEVEwR5sA6e3BpdjGVBv4Z4oSN11SC7T7bfqnssFTxMC
sFmxeZvBgRGgFbKAI6wFhk00jjLgrmR5ROaAMUDUIUc1Eiv8GVqIFY1UnM+k6y4g6rHGfn9tgEMo
1sNmjLy7IWAhD3KC/hKOPlFVHnIjhD9o8SzCpaSipL18TzXSFehaFZqdlash7aXt2gjmtG53yT7N
2QXZUhpB2NfcG/Jxy8egF/n4/AdRVaTHgENKEg7nZim3uxmH3i9WpuNhTHsRysel0w8YEkw5Hb78
FgaUsEFjwPbSXbb/RcPjqTTl8L+G96HBjmN9jPcsdDwUDZ8SNyLTvJhWJ1TuMJOqiRtMMDP/hQeY
eVBLSwZVfiT0DT+XSqlVT3lTaI+cmm7gLhNkLRrXFkFJHgzeltNWBWcI0lmrVNHQim+YxlnXYfmw
AMIDy2vJTyahU64yYqSEPQuDuxn5omVfETUrSLHuQWVTX2LhNJI36SoHKObGP7vngJKT8bSdGThp
WVaeFJ+AZImhEYdsGYrG8SwHvaC9HW/X1rUA2YS9P8DON8v6G3zfiFXPdT4wfdQGbKnHrP02JpCi
IVB6qk/ASuQEMg1hH0snW5iObBgumSprdOiZI4X+RhDBGB0ADn0L8oIDbe2xmRZUia4raAKFheKD
deuXuxcf38sv78M7e3tzaoVosKcG+TWRk06xTr1v5FPGaOlvftnE3nq2O4MA3Doo9P+u58Tefn94
cSkySAUUMcWwB3ks7j8jDe3b8K+Dj6ezIKsMBYo+Wx+uwS/JsftiSvZu3XB2dFcztcbyXzA7w17e
C1XhMlqRCI8M4mJxkKW7f/mgSFTCLRjFQ1VfDuMz3g9nd+8VOmddQAh3MH758VzoZj3fZvWPmhzp
NxgBZ0SYFcX9Nmbnxi64Garvj/kBZb/G8WSV1fBaY/VtR+sryeNpdt5TWr3EqrNwPkmzNuO7wJ52
nlFfPWvTCewogs/StedG1CGa+TVuT3hAYeyJz2kgDbhO0P075ektTwXi5k4DZQ61ZABtj6zAUAfr
dxSDwo+QXP4I1LCHk6USlnO5Lj0vp6NVBu0CsY+3Xjzh2cnRl5D5Oy510+msaJnh4+GaaLRBIdQe
SaWUajffJaIQEiqGq31/eVT8dp+Yvo+cwCQyPV7d8lkrWJJqN7wZ0Qk8y+TmVgamQn77ANJk+8Ld
iwHIHB7VcmcGDkCDhTeFgdQG9/gKqzq+3njXSE0cW0ooAur5HDwCML6dDmSXQXHDVf5N2elIIgu3
GvEM2SqYKHNmaAvcyKQm62RZHG2sDLQ99n59VDMLluxJGy78VnjJ/6iZSk42dV9ZjcoreYMMUyeV
jdHmazG0gHRSjDd5nHLUS0WNpPfGQkdHzmrWC7xDlZGEtrA5UmY96lG5CfilkGtisxkxR+xER1ov
mvEWVlCDj3EVO9UMZGx6cGYwgrNILFo/Ix345klAPrMj2AE3XuErIP+9S1O+J1xBVLk6blqGeOa3
ieOuVrmVsGo2d8808DqcGs1xkr52vQuZo4Fr/Rg63p1zpPQXE5Nid/xMs60EjglOVFc7cLE/efar
boT1BICRIo1LwjX/LwKrJ3QWXp7IWUDXa57Lc7aa4muu2s99RFMNA9nWJR/k4gYeJjg6LKh3Qxj0
UgXQYJ/0VvT9uoMTOJ3KQGEb24IsDC5gNhwB7fnZCFg4kuwVg1HEHaAEuita9viRBbYlpiRvTrNZ
93TPb5aicT8jvEDdrziVQm/etoDU3s2G7mwgMVoGDoyG/c0pCeNQHPRopJaNKgWlQhjKEu3R0FGU
oIBjl4qvuLeuExr9rOyGNrdQkeoNzEL699oNowN5L1w6f/O2LfacXyDKcmqggVqCSI4gTreEqC7o
RHt3HpXH3/9Oxo1sGTbH+dUHaEtZU2Z9x56CYZ6FC/MIgw6PTmJmOS5qiTE5uY+qJSC/GLFD2Dcu
ALEwPMqq/vEKybstVGuu8dHqe1WaFm7htgQ4/LLS+BHhPiUr+f/OxdoU1NWAZFE3R9XZ8bzcLq3J
AjwrlKmns4hKocLDNjThUOGOn2BJq5qlj4SJ9HRUW188DSqeNsEgC1vHsaAzffd8nZUVQZBK52Zs
HNHtGnTKI1CIJxm+4IhJ4+voF5Exf5g7ypE90iR9B4qq/AiN/x1LKJOtCk8gYJgx8Kb2qZb+E3Qc
8X1fZqg4ewuYnNya1SeIwdwacqqVSh/3Gc/7U9rgC0y+ZJVbffyPElzOm6mVZj8uRfaSfkgw8Hwf
OpwjA47v7ISKyVRXEbGhJMF4ArgIAVJoVtrUqVEju7nJk00NQfMwIAf98ot8oZ7WncohBIQHZ3jh
TGGzHKWB27QFVT7Kjm26j15wY2jbWxtJDsrVyqdZUl245whBhbcklKAJNwxYQx5tauVFeXW5miP1
QL7n+SND+aoyYzXd8wAg0v9CqffbDCwW0FuOH1molWSY7fSA/4Z75Bm2XLLet7hWj2LLDRgOqxNk
NatJHmLd1DVw+IYtx9uHrabMak9Gtrlnewt1+AuIKiJCT/iuoeyB4Ruebp74MuqalZpluAG2gq5G
A+NS9GP3sq5mDMiSQYFkYAjDU7dAgqc0x1yjRnak0DVUmiRfeseMAYM2pfh5tQtfpaXpRYR0tw4Y
2bNIP7/gxs5gxSSG80oiZo+kCgLvflhLs8wdxi8MKZ5LFqUmwoz3pEw/lnJB9n/jxtOoU9xksZgp
6lG53Z7wfkYzp7vAMPRlahbTEvLB1J+YzWRoQk1CM/1g61/uFKwbbKdJLx47NySsY8YJl2RSIOnM
xag2pzhdQoBtISEm3EpSq7RB6S5Opj8g4UImJ8C6yuZjVRWVRns14jAilpU5KJglNQ5Oz+82WbxJ
nLcFTqcNZz/Jbyg08RBsIQoA1UpXXUD+DRH8N+yaZxSDlvkOVdZVKBX/HiTMmvn2YEug6K9NMUE1
P5IqmR8+Bkz+Z/2Yj0UFcgfHJuVoiGmr82ykhW8xNQ8DiS/hKTdNupQkUlM0o1SwRxmCev7Or76y
3yH6I/5oNY34rsxWpzghhF1LCXiAA+c/mwuqjXUEF9S4sdcgwMt99s+yeN/gISfKVKLn/O4D40Bo
LNZO9ncQFbGHbY9RoHcmVgp2tn11x4Ij8NOS0amjIQcGt9+dcB7upK66OwyfNjSEWGZfR19mhriH
9ZfXPDa0PRef7zTqpzfD5YLRvDvRWIvhX8MESFvYHBblg/3pDrYVHjVM6nI7OY5aEGpDGyqQQZ+t
lGwzMDzjAhpnckG7rPlje/3DXHWnTt5pJ3eYr3QMhrOuf6HMjIV1rby31eEiMZzOb11udAh4LXm5
HRPV0X+FOaFDkU4aG4jZt8v4ukGKXVOqW9v8QWnAbvAN0YSZ2XOXOEQVpAQyoKdWp6swwImDICZY
alfCg2v+0iVIMn6wPtXpvs8kZ+9s5Ku8o5os1v+HbLzBKQ25f8uN43XssIXigY49D3Fl1lWYuQKq
Hu5Uzsq3p/JYTiS6C3604nhPmLSBjzxMmnPHhnfFiL3Le5dmifyLSUcl5rWu8Lo16nM9EYjBH/sw
VINemGBi7XepkpHO8KXeRbKSQeBB9AzjKO3NVnuqQLHRAbSkgZZmPiF5R6PtdOu9+Fq90dKlsWaC
6vx1t6OhWZbNPBWX3gkgdBtid8IyNnaCvLC+gjR9ZNVwSkdvxjX1k1SLtwpMUr7JjhMKKf2pALdh
de+1QFidfk1Ejb1UwNVzf94FkHY9TnTasjj2/eSdzBN4tej62UV6pbEC4FsfP+JIwIQVgo93juGs
LpDMbSCYpBQsocZ9C3vE0xjhOgTrcs+ZnkEwoo9xf8QOS9D5iIhwGssdspyppXbis5mEjkP67h5s
xV5/5v84wIVezdnRhzj5MquTJSqe2hmz18tbC2eEag/uVj/+qtVUa560jhmCOspco6brvZ7pipWA
mypb7j6f9MV5VZyPlkpaDy79t9hNGOhkWJlG5fWGjrSRTESurv+5BI/gQtn2wgDCSdWXzknBlQQT
x3fe2mKwRAIkydcbaFeXhwHS6VhSg5Q2CXFLSHZTdO+m3qsWvkT6izHJa9NPvhGBErUidCIQVmxt
ealMSx7ML1LdIWYYV3VQJgIKZigi9rqKkmsOpxvH7awkgcSQwNBn3Lmt7ZhiW5PyryBwDWJ0yV3e
EFnzOhcXvl+7BGxrv+byzdhXwrqVUSBBZznO2q5yQC72zrmQ1Ye1ybsoKuKGWFzfe4459AMF+IJ+
TWGSsac+1PhrlflDQOOMWnXjy2P6RwicDNODSWRnZKOhP1qGBqRhgUeiTHFzOXAdyCIPQuIzRG3R
aDmovJwx6Vws4rZjop1WOYKMhbT0VfXzRmIuOMJw28W00hPd7M1uS7+WCBX4/hHZHXAywbSbBMrn
yump9/Wyo2UEg+5kl7kHJrESxnLsD5mnN0l31kLizBxXqdFUM0dxEu34SHvlu6P1VN7dqZKMIL+C
DHNFam06knmpE3lJWA2ThRQTxuit/fQ9M+3Rg1F1MkXDQGurOyICw3CHxlEycd6cqaKh5NehECMT
EhspTTO9b8Q/qSHgcCH9ZSA7ntiXaGYyvJZ7eFopKOwkwPrP7FAixKkGMQcFf+LN+Rtupcrr2cCj
ykEowpQphOBLG6Hci3wZRSjKDbCLYqCelMbscun+42YB3WMO4D3QvG/E/y8A6pygr9Gmclv+UezQ
W7w3icgn0ldgWwTtHHjf+QD0f/Wjvn+mWm5IHqRmSeAfDb23MBp1kvM4fMcPx8S2D64LBDBqdb7k
1Q/RfvLz+5yl9c5sO31tNkQG1nfCbdc5VT7Fp1SmgT6+0g5n/Rf2qGBSninTkAiBIGBrk5kw5OD7
hEgRQbc2EhRmKrBl6R0EpWhbiPtRvJt1I+LMOUhscnqb1aJUkFAU03cCIBLJLjwW1vmxiqOAav9g
ZEYzU2DXMX3rnroKsh+k8eOaOcwmRT6xm9tXc8hkdaWW2G2SBBd4mzbju1qAomWPoprqorEJ0xkw
5+9yr336nPLEsnD6VX6E5CMpR8R0yOGC+9TTRDl/Y8u4S7PomjmiKlPhxj8V3EWgEDLnbsIZ4di8
Va6kHMSaUutZb5ern7q/pjVRwRFWeukQYDqPwqjYjwcbn+Pqhg7Rh3i9cb9OR/dtm6HtJo17UKs5
mRmVOVTQ4EwIpG9gmYjY//+xlCJFASv2rXryVWXR8bH+Sb11WpW/G8y/p/3RAzcrRiVxoIflPuNV
kK9qEb/essNol2laZNtFeYDHCd2gX0L/dA+WRoPKAc/fZZoVd2plwMGds0yhf5t2Y/5sBVirFpHr
TCpCvYofS9KXInMEEW6iwISaoB7C7+dMza+cTWbaR28nhwmEYnAvkx0/3r6fA5u8UN4XCzYy24Qg
z+4ZK1BAXSCkZzMtpwTNjbPbHCX+pvKp9+zTfvuzNZgJYTz5pjej+LXjcSPOqB7/ENmGxrRLmhjA
8QHsiqeviSUbAnmsTE2QVM8mpDGrB2PBouNYpBDAACuDvdg8sCQXItlYmpCHYBG7BczmAYZk/thy
hR4yZ7HsvcwgGvPvhZ+tns8FrAEXjDkpyZNAbjyBPMAoZaeYa2ZVRKcxHWsxlAm0YSkcI+RfEeRe
zxWvKq5/YC8rwPPCDS88/nqp587VNs8TFyjsBbG2/g4veYnBdYxhk6p0AsyRBLMMPQTVBjY6P7yR
h/W7cJu8RjMdAvkk7u3OJhwqFdSeJk59+UM2/QYq6VCdAEHU9oW/T4ROv6OTuq5BcCKdkxphSrGO
b0+/geVCOIEdpol7j4eD09f2c+gMylYFsCd6MAPdR3sOenvFh9RIJwIukJTVMz3cOvEMGAI5qIKv
mJI/Vzw/fzwvh4RJF7zIhG2zWmRTYQ92c5+q4MzL2Gv8g6Sdik5zBuIuuzmKgckjrBjg+28NKVoC
LEdGv/CctYOQD8IDgDyD1eo2NTCGLz1UwaKoNgOktQJ4bdsP4fLEH158LXSIdQbxOb5/+4NRtQyX
bXgKO9TwPoHqq3pgPG3JjOe2EtR24SnWPxsFWECrN7RCuVD0j/ukRTu0dI691JjBUjs3pb55KCM7
FIPD8KFsOuKOKzQxvCYlsqT//U9gwltZmez8NyLHwvkZJdPt9h7wb6o8oxQFiaX5IhYo91NSMLWJ
VlGkY/G9anORgX/vSr685jvpgGXfLVx8dSN2MtCfvbkdMoWkrI+G3n1IDlrVt9sMI0xOEMmlt2LX
45MXwoaBzNN2rO505tGn7C5EVg5Ekyb4ZX9epjzB5kxsuToleEcHvmezOSXSVT18d5aenSQqXC5n
W8DjA5sXR4V6ENTWU3pAvEt4YdZ8A2YG6DldW95PMrSnqNrCtXvjj9f2odcqi0vrgC3cp7zn7j3p
Yah6tiwRg5UbTC6Yg5eo/EFqsMekDt1VQGn7cMFp2KkmqPt4YuRIhBigBzQGd205TShSJ+r6MLUT
JhPkmAYdINbtbs3ADwo5Hjq+FeaaA4McF0ZQ+StNOeHNnVwKYBxC5pJeoqcNkCRHc3ehkno/7GSt
qL48hFSZFpYn0YkPpSETNn7G5fyOsZHY1P/ZgyiIyDvupjP4PHBqGC36xyojw6CBa3grLydewnEx
16WZcv3lVDJmXoIL3+j9XoifPmfUppKXzyuqhYk9w8J6BAHJ20PzWXa9DKu4QJa2eoCay+7PsQfs
7ZOfcHiyb9EJ7J1EQYfmuSnA/XyGQePGWKqTImCUiR+hAtHGNUEaZOwG3ECaL8Ru8S2pHC/GEgbl
91jumzQp0KQV9shMeWFLMmv8lo+J5mhDhBHUTosez5JRqeAgosE5EknpIBRRE5JhiGwIZONvCf1B
prybeWWljmq2HHHn87JyiNwiem3ohQgQ0zYOTnrqEcQvLE6CZAn3XE5Ts/Z4zX2mcyDupe9H2PHJ
niOinQeEMDQHNCEblmNbgAICyd8gxBIKD2g3xveIA1DIUJwVnG+nlIiN8XCh4IaLWMsBzEwS4Zqg
Bv3h/T8ZwX8K/kxR/wIcSSSGvIr553jgctPIjyFvK8rhABCQIZ7keVnJtPlBju5q2JkxTR53Eq2z
oQhM6durJEdqscEIk/DhL4v3saUic6aMM/J+MJ7lh0ycgygIipSC67LqgIx5oavpMmccKaqa+mU0
+SasSn7VPtuMI24kJJF8gRPD9Nm6yqQM01ObYPAMfMNpzBaw5xt5Y7WIb9KgjTgPBvv/MJuLFvxj
CrjD9QFLZUXggRfGiTc9bT2x1vqHIGFmH0Yi8NbBG+JYPceYyiibGULADnYkoXpIVd9oNLojUazA
DVjEUjeuY+VSWndY98VNm+/oaPhbRQ2fz6H57JHlLktxTIVYCHnk+mhMIaMF2LmFWLcFaOraq2wR
CktnLZXOg/fogzeWcNh7XvvU/jSF/sxqa8DP72nQNFtsD5APPcEpJPJTkxpgLR6264KSaBOrcBLn
l88E3MffJ5IrMdbiScEM42i46Eit2N3pwuObOfa4ZtfT+m/xCgSVcmtAI2vuwYwz1Kxt9qlbtpxl
w8RHaALLWvqKeOqrnNV8rplg3K+RCSmIHfPtvGS1faFLQbId3BVu8rLe5jJ5BygS5rgq1JGtF/3V
HzCzkzvnS/BfUIxBGEbDnMPlN2pYpyeJ8W14b4xO31mVH8TkyBueKDfyUQYJ49l1pU2oNmZsfjdP
1QyAPBGc/u2fHmLJIZcOEZnXHqheRXd8jDkxdqlKthg5ODhqIFfHHNET2gafczlfpTQRZB9Q9Kl6
MWFp6VYcrTEK78p0wrM9lJxMv+c5pwwI3fugbBSBT5ymm+6DvyDE/Sv2RFpKns1ghbLztowUei2S
sjAbJcFe3vrlterZl2h5DMTFlgXt0nxnWhsYYUbIECUIr3Eot6RF8GpdO+MPaEJ0FZb9eFAHp+My
W/+3HkWVWLOG+STnbJIoSVNnqQYVTA7ADquFFOFLPyOmYrC9cEN5jEzFaObqYgw4KZ7az+OptXqb
lNBg1MSHpw8WF+sVlB32TbE3JazXMtWWZ+eJhnknJEzEFaL+kgWsRXRbdXgoHgjHoqtpeMdCrAlD
m6cV0vDvK8nbWKnt4txKjO+z/CfsTMQQNdSYgfhd5m/oN4debNFpZ14fGI9ZKMscJBNBniMxzxxo
R3ogG/po+Aoang30mC4Owf8cmKb0Wmv9nKf+9adWgGaBj4zP5AV9GWmm9iHRMGWxnTxhrO1CWMRz
bYNOgR/ZdWq1eQ2gNQ+SciXXLn1E1pEpRV+BTrYLJL4gyhD/ghpNT0uOo7YYbsnmiAHpsxioovjv
zSl7lv8Vmr6zCCQjtlWXG6qflZqvT1GBrmCNFFSjSjY99VqJTXCZFmkfCSMr7687eBPD2qyaxk9s
o9tW1FmPBIZwOujt/9XoBK56HQT7FoN63LuX1xyE18F4ObwopUlFY63BPnP/5aqJP/GZD/DtikOV
GdYWHVdskoTfSV7+U59SRW9AQoPwbnvGulbuWXo68I11Y7W6fQa4Z89HYki/H5PZ9vtnPhQ9/aQQ
DMtNxVhHiJ7ugYUBDwVBeeCLqUVUXgLix+qPV04r16thRt8ArV+lNHtA9cnMrggx0HwLnfSD/FN4
wV7IzKylChmYZoLDmkKr2RH3EJxNHkakeSk0QgR5eCEVa6OoyGv9ggs0blG77CigDF8bT8+QLzHt
J9LWYOR4q+Ov/D6O4o9nKGrcqGtc4ARfboGJRtAfV8oluEif4FdflCGj/qXLR5bSI+DyBnCFLkPx
h2fwWvv4OijknrR6TK7tNzIvpfnLWIPbTN/D05EjqwWy7mTVwjk9OMbu/xHNuGbWBqGHOGKNgJtH
M7KvH+NOpYcZ2KZ/lJCvqNh5zhw4lctLn63Wtnk+Jlx23cBOnJgVoExB+Joos4WUxQdOoBntjrph
HUrvCTAuQqaLHaR5t6Ib10lMYD1ZvgXbwr1vww4O9HbjkX/8ckxnvdHnoGDaNc7kzj3edPBaOvqu
CnBN9btbhTm8SEt9mPnzMDBgL6XtCGpEu3Hsv7MfcWPW7rsN7t23SzIaSNTZnoRfllkaFzLvUM2/
nbEUk2YoTqOeTd84KKGcX/gesjp/SCNvWFeURxq9UhQt29/k3rCrbqmxert9qV8qH56fjaPBVr/3
TNMWxrqhwdZj4iEtccrFajp6Qg8g4T6td0W+/ok9ZuU673ojD7FW5KbxKXNBy+wfYpm1W3zH/YXi
6GtlaPQmYfwZM4Gzt54sY0gswF4Ggr/4/Yds/cX8S8SNa+PMDH0QA6WBpjElUslY2kkpMrojnHnL
05eXzvrNAcDTK4wJ8wEd+2rPH5ogjU6qEHQKlbE89m/ue2tWST4g/U8uQ7KrcA2nXBxBXmRpvWa5
+qKCk02/MTIuWyzriKrID57bHRoXV+BpPXLlUDcphuczsvHf+Ocfyloa2LLHhKMaq9bIiB3mruJj
Yj9AhbQo0FCHRFVf/9oGPJZTAT4Ek4LpRZryh5t7i96da75X+aVNgkxzPXfQNGZjuhbzIrmdUhlw
7D76KPxqaxrGFLYMVXyl3RTt6bTuP+N8qyI0KCzIg2VwJOglGf+dHYcFudGH2IywcdeCJ0NjFggE
xGRW+99nfRKcfesVps9DMVB50YHBzaTkLTiZFMRfnaGZgCuX1qHfQBXhzTePqKmYwSGFId1bJlYw
utFTm5cxIotPAlq5qPRG0nLPJVMKSEDI1tfD5//62AHBuigL0lq/LkZqcfOu7hmvbzRY7wuywsN+
wvEtLj/re1d3fHUmdEocex2oqD5DqBRZYpavcrBLvWyJQFImAYB5Mp22lUcDQzUV5kym19cuW4/T
DHkA9GNDB6VW+9+Spa3DROe3CSAZLoUShtsaNpEL4vM9sRbQJLEmlL2InQMiLhHc9qaKGq/b/4aY
LlmGTUeC7NPXm+KP6pScefWwSMd7nC1vHBMQXbUmTWpDk30ifmLoVsIghdDlsOaY/XauwcmCELJV
nt6Y7Z7o5agwl+I2NzmySf8ZghX8oBl3qUrYREoPk+GUYHPuTYU0JAxpjuOZhQiJopQlxr1yIFH4
ATHpetQxNx0o6Q+NQGx5zC+s6ehkFT0c2pWu33x5z+ji6+RFmLIru3yz7exJyeZ/3TACKMeutK/E
CTe9tfYMJ5mRI/Qx+ulA/qsz6grRp6AbHqNdjpgDhN7HTVlrTqMLbGas9JFqh26TA6zHNvKY91Gd
jtHHkgT4K2nA7GcKiaDb8r4Oi42BYMAs3QDHsTOevylsrA0lp+dlYCld8ulw4SygkMIARiwYkV0x
6j4Sfttxe2dGTIUdJOKyYpoFCY6ffzD8C62g9TiK2ZJTfYDNLDsYtn5twPYkirw/pR7SpXa5S0u8
jexDGg2ItfVYglzgrfn0SHAf6GYBtgsk99i0KlYfFpBORnA81QIJ+bZzprFj2HdAYKe/d/q2fvnX
EGvuNN4hpOUIMi4EAVfzxmkg4EiCpg6Nf53Hp3LQF6MZw3u4to/H3BnP0Sa/vHxc9o+u+ENMY9wT
MDJ9Il24cw6Z8kjLFnSSxEbvubpf6t/KFDt3sT1ywLrX9IQO8AiLuVp8KRi2cGstfyD4K9BfhnX2
YbjWUMIJ97dR+ZxLeKW9UqpAtjt0NC8vz6VkO15HtxLg8e9uHihQxJPA1gO8DPU6Z8Yz4tiIE4gn
BNNo0PMuRV1ozZHfH7aYyr+xsws24l3YyEYQIwmJbc3J3dBW3R7StwOc4AumDwkpQcUMkCDxnYwY
pBEALTWpkk5rh6+pLZRfTd5Z6N07Q++SZNzcPVGRBB7htF+pBXFI7Mj7HEvkkePyj19LBZwMYXjJ
m3zFmeSGxcb37IUdyVDj1+0R3YeAAn6eIZa+RE6DPLYfoXu5IIl0K6kg6GpXHkHAvr2JRQgAibeO
wr7W+bsNqh1OUUUpMpkeTgHvTvMoaIOMiVKtu89OD14LDBacJxSxz2TmUBLmPEqttrNd0h9yjZu7
eqCgmjwLEaR6RjLw5fd+xUpYcc9WB4GkEW0w0liW8CxOeWUb8whD3iWk0vTOIo2TB+A30In2+pDz
D+7utKIWgaX8DCc1k97bwMpMahgEgqHBiVUWTAAZ2UxOlJqzPp4dTNOLX4aE+P3Fu0CeMLg0nuss
Un1Vm9+v12LQTEVvv930/FkQV/Q8Ih6H6N3mnTG1AGsMav6H0iXXAeet05raRlRdYbgz5CiXgJiz
IKWCq9he/IBvYq0t3Pj8M/Drx2CS/1llY2Q0tabMW1L4TuohjlcevssxX9S7g78M5RBG6s4NyaX6
o2+mPkxusnSUDybLILhDoPhLLsHSznOOBazj6hJocKAj9xncYbfIOMWVjPr4isMEFvvaiiGeGGZe
kxvedcGluzW+FOKvD3muGL+j7kByL6T4sv01qfw+d1Jg0yt/ZxH0bXENjOLzr396KJVYbgT04UDV
hKHjhjUQ0Mbh+XJ1W44F0C0qP6FRE4Z2aX5CNCNKHih4PZbmSSzr7w/oUTuawxyJtIN5A2oIQtEj
3TWi1GyGVaFLIDTfEybiRWpTetfQPdqSmG9137xAgMhdsbFNsOVUVNK6XhYzcz9agZuXhKbwDyMz
RhAXuB+h5gDDkdTR62O33IgWEuf6U5n2fXSkAYf4tXSyPiVBcVWNAMtsrFxo1Oyv2bE6/76iPvjP
v5fnj9Dx7ZfS4Cw6vg/eIwBOxOXv2+Wk93gz/R0yRXL17XraZfO3SOFRJH8H0KvPjMJFYS6tPf/C
coVU90GzZ+r4cwkOgoV4h4K9/0fRzcJZQ0EpLg+mTzP/HwkIkMlNVH244e9qKY3AwxP2IVpafsS2
2GhMExJ55rsFrY3QKKkdvGnO1/hJFjyaxHN7xeaB9T3f4bptcsCmPn43phCSkXZqMwlMz7aN8l04
cZkNoFyn+nt9KAQ3+ZkUGk9h0Vd0Vi9Ov8sVcGUQaoNi92UM3aR6ALkNZxjW8OZCaMJTfE25hcJ1
1ajutzCikK4Vem7k8nVp62UQURGKsosEM9M4CeYxdm6KAmhCc6+6L+rF+9IaoHdz1zXgZ9iVhS0Y
l118mQWqVSX1xGaPCrAaKrfW6AYh5NGpNy+m613fb8Ji0f9vnUJO69MjmAnKFwFwf05gKvhafosS
r2WldgQsWy/nMwl3/skIPE/sFESYidjofGWs1/WW3wH5NzKzPvmLk4lwnyka7G526kVdGakafO43
Qfy9ed+/YTdEOetp/PoJQ0AiWJkIRYJBExB57pFPB+20Sqvhr1apCJS7jhRL5fapbPjS2fcLY/Mp
HtWx5zd6L7hp1Xp+1nXtlgSrtFGadB3zQ43ZnXIIIngy0FxsBaONX6cxahrcMW/0ttGn9SlXv0hU
YGGM7kZSBo0Tth24xEs8+zNrZKwwsLj9UPV6xLTiXkyHcn/fAHhSnXW1v3eafI+vF6oMYahyaFY1
QSfeKLh7w1/5KMcnSLvs6NABP5Sji93FLF2NM7d8uUj5cBwthJ+r6Q0V3RecyjUXGDCZYcIJsBYW
Hr61ohUwL9LmXBQpN46UUcxe3ewZ20XxDa+tu/3yV1CV3mC8Vghc1jIWDPtBhEcLKUnlk8S+enX5
+XsojGrAwWwcX+lxA3ZnE3W/WI9gHxTqaL5dPepKPuTOg+zDyUKXp3paWlxsV2fl8Goietro0fEi
o/r6lsSkEUfu8khdvJ5dg/RDr7GyalW6TOS6Hg9M73plPfe9V0ylz4xdyCI4pQSoSOK/lx9T9ajR
3wdzubAOuPsIUsDb+/8xnEsNmfNxYXIiLlmgVYFJXhlhZNxxO3d+HjNst11c+BPjwrfWD24blRgH
ccAD5r/BWk8NjcNPbWXVgoQc4Kz46j3fjXRGwCm59R1CaxnByMrIm/kX/EMNprrV2Ht0l8+jnm0R
Bh0jacU2llSvCw8nWzhS3+d6sdlTnL3w4cK/nm8hRtvCWKQ7yNYQIc+ZYt6VqVfN/z5jl47zBotg
pnmPVHuGX2JiCtp0uC86F3CVPgM0I+lJOZg6+4759l311P7c1rCCbkUw5/PW4MqUvsyaQQKZY3fD
SxWFQ8/c8J2LKCiWY2OhH55QADJgcIZGHbXQg0X9DEWHxh0T/4iHOCMuhy2t8y9AgDBQf/eyyBGU
3kjPo4kTkwztIjxeMD9ArCRLWAtNk+WccP1AWk0qsgylJqL2A197j2h81p/CvOh9rdjjjuMCnJRJ
yQkeXYnFSd3Gil1cH/tY7UFFZfl9AzpoHq+FdQ7FjXABMlPeQucw8S8o/YVF38Uh+SfyUsawj0NJ
Vz9s91frlvpp2oaFBGpPsOkATzi/R/U+QfaIjWnpyldOsiMfVTyjOEPVqTjF0v1d64z8GizbaeRH
c2hmQmrq4+vrDPvvo2zG6EkXnl7jJViZlrDLDKttW40xGkMMl6l08tUBzUY16xlhapwt7oFg01/W
UJaX8YPC99CDNbKeGV75VMD4R/hezQeHw4L9wt+bCmD6xnfjlxsGaM1L5RiSJ78LYMWLwaKnAaN+
hh9ualOeDjWMjN+rWPUK01uISfYHr9AKkwbNNNXBDlHAaaYW5WkzZ1iwUXlq71Q96UPzPZGCEcve
6JDxrSWxi5uygEJDG47DJCjhbX8h2GpfHUmsUE1oD2MtJLEPvKBZr1qcqfdDV0OhTuMy/1loMB36
ys/CcUUxzMEQh0BWJyV0EA3Uu6FciOxNvpj0URo1JB2bRbw+SknRJL1ApFVqRap7fy+gi63glBRu
kYII2Kmbk3vyl9gOlAK6qSxz2TVWVIDB5aNFMczZpVW/IM3d7KAPHp+2nyaYeC00FvlKx7JtL03o
xHo9yLnk40PaeqQrY8rEkMR5f+JaO0RtuhDu9NdbC+B26G1Fx6LD+959ORfC2JsWPqIkL0s219Kw
bzWjjioyR66VogolNqHs7DiKUzzlNpBeEmWyaG+ExepWV1LJpS5799zZKstRsEYktitGEvpN8a+Z
v1RSkBvDP/HSCTeHSyTL/wkyrpFnXChu7QFBet6OM6L5/s+Ife5s7hJDGwr4FpW+HBSUwAAx4Hzc
wuMl5/ZAEp/L6MzH9rD+E5LiVG8WynJB7jMaF0EdFrOUzBCz0ru7lBakFQy5GUNDMep/GwbLxY3f
uwJOuZnJLG8ropn904kfnNS6N6tVtZdT3IT7i1DG3C8BjPAje7EKhqmA19hz0anu+jx35HA2tWjt
Q+ErADKD7Kne+5AmYpvyISaKVjfssjopGdbDfhu3yzA8k3AfqdhhQlgZFx/3jdeO6oIbpVOO3l7n
ann9UVqXORDbOIa3qVc6v4pubBA4CJtiNH5GvVwZ27FwzNqIjHl+egcmX75liTOHhCnbOVhT9nPe
lraw+Uez5k6AjV9R3I/VH+0hSt7DIBz6mE5y6+nc1DNhQwAC/XHKtplGAZDAJ+5RmgxxUyRuE7Ex
B5mj9OO8E39zqU0KaIC71/pvJJIm14eYrwSMvrFsrG1bAoQisq4Klrtj6qoPfuCaCgTOE0TIRa0P
16ykON4G9VEwm/5NkIktNAHzjx1pJNq7YlBdisgOpRFT7hgvEYPvmUUl2Zzo2ETqWgoTVynZj0+h
18ei/Ovfp3iXSYf82tf21QNPPZDHJu1zdnGinuoyKMR59GwlCcf9NPS8OfVMKUv7le7Pmrr9NFEa
TCYRyzqthqOxTkwZEf7As3YI9AGWCLvs9kNpmMB5lCDFEABCdpZo/hYuCdmPeWp8Sx5a6wYTn4Sm
bNBteVXZoylFB6PFmBK2Zvo9BSzYu7TdJFVr/RIYcpaoQbn96SQkg/+gB59/Q1ZGD17d+ucSUVno
SCv4FuPvX41D5foxUWweHbnpKTWpL+etJlaPfau68HgBqcIMn+lFFyMxnDQxMY/2eyBEYwjhnEzF
7QwIkKeovVrYMbitmgtGtwwZcNzemdnMqjZOrBE+pgyqJ3cYNzg9sT4Dz++RYZ0v0pA9tNqsAebH
yW2p927uwdka9wOR1IVQlK148p66JqmuaXBQqm4nzTcl8RZTybkt5M3B3ZkUJt1pwtgB7s7Fl3Dt
85hx3hNr52IYqC5L4KRNiNDn39lYs7qkucQcGJquu8O23+BKCYqrh+AKvJjE0+Nr1ia3nyuHTmNc
Nlc0xXfVJ9y/2MzQL4od65tvrwCKtN2bFEDx3e5xMdZd801i9PSLPMMUPZbvHMRtSoT1B5RE+zRn
GwV/S/Dndat3HZo4h/BbcujDY53UoXl55CNWFaThC3D7zOVBpsrr5VrBmhhuUGw/DRCM0/4fLd7d
iXCiMLGcrp8JPW95asaIbVTnZRKpoDPnbY617tzE31RvghZje5tFa28Rvh2NmlsoMdui35hO13be
nlIA1ByS3uh4etmV/1ONxxqPQfNn67F2x4Zy17IxPgW8L3wXVd88ZI7BMcCiQQmmefKV3plr87Ke
VNKHtkcjy95tX7O+hnRfI3osQo87basVsBGMdeF6Qr2dfQxzD/WitZxnqeA/nsQ+l9imphEy1Ty+
aoYL+T/lyqCo6ciXEmFaMu20K63pJIe6Eb0ozsp5BosFHhQsaDFaCFAunQp75MO1N6/NgnrV3Gbd
psKolUaWzt9jPOsThlD1bRrB0taPKQyBsgM63ay2HC3mQZQtPLK/FbhUFDhc4Q265qM7SamI1g7X
tL3hokCs5xf0eKjgYijE1dnGJnypIMjV7BwxCA5/w5L3c/Os2jEckUJiXT+hmJoXqI6g/CqfjM+/
jiuDYlzQuzQk7Bugj9Jw82rmxkJXX6UyqECrfu/ssLf5M3NxPSEKgo/EWwqoSWFdQ4ZcerFt2nr5
CyR9RFWT7xogHUGikRcs6f+j7a004Sv9NWIJfQyipXK95UIw+45V5o/pIXP1m0esabRMBy0sR/1J
e22Bho4HmV1s1QOKt+7tcEQG+I00jtUgr9Ng+VG7ZXyl2cU8Q9j4DmA/2VZa0kDNONo9T5SQCjrw
R8uLqkfnmoNobLZnm3azpsMxpL7rQEUIiGwM0/R/XPbExWGXzyGkejVdZR0TCU7WmnTeBEW4mqGY
7w0uvDEdVil2EF7NUgLp9cjp1+tE4OksPNVvdjBgZC1ZOLQkYs0PHGX7rsuK7qpRukXJx/Xnnvdi
Ik6Ej0xwpa80PH4mfa8zZDYHuqaI72G3ULcd+cGs/01yaAsqSgiwR6AdLhss3M+i9UDgNZJshZ6R
rgUdPvf2EETzitjcl9HCaXoCs4M8HdGsuSkxK+TkM8TyMRg9WbQxq/j/5SeKQkhNQjlgCSY2yv3P
y9MFGiLmUTWwIypHlRgXaxn8zYeu522fQRHU3hGfWesxkZ0wxnLT0UhhDHgS17kQCSYHDQ6e+fa/
WjqLxYEKIIfIFTJ34+YF6Mzz1WYpaCT5IkE3U5rbSxUH1ubDtl7+fSJxo3W7LGdypEzPK+JxzRf6
qTHKgUI+t8SpaZzoyOo7Ba+dofJxa5nOZN/bhU3oGDMgI/j1HejqzNfy55Jm17yJ0/SD/tbzo8wu
WW8m8xsxiCgzU+wiGT0XqatzsmmKWF6/8UnucYZ5VhHUrB/f4eju0wA6ja2+Ughm3Y/5w0xcUCOL
MKZkNsoYsWMJxUvd/izQPUBaXwcEc1c/VU0fCOkGXLoizyaGIZ/tp55ArAUkCF6VrNPxB8LI8fM6
On1kZ0ppj0n2yqV8fSl/dcuzjip9JULNhreEebs661tQP2iV2Ks86jtzpKh7vZMSRMniRhj0Eqwc
EV0c8rp/PLPLulEh+oGEJfnx3edHtV10kRRHpQ0meSgpjdtNile9YBQS7Vkwa2ojzCkJw3CSAPMH
tX4jYJq+I5A76Ff1PWCdDE6JD3/vj8OXkfYmxvZYBALB34kCYN/7rjfNadcl3wtB06TtPlsbqxNO
IbgB426ey0vSXCzmWeqw6XtCEAHoIQRU+cQcBx/BENWO+Nbhene902FLGZ/ydbPMft4/49J21tJd
h4BggbBVn+Q9TVQ2Kb1pI0BSCBgwYCWepmRRZFNNPtdsjl57IXWRMq+VmbTKsYCw+MRBw6XgFIcQ
Qa1EHgMDiFcRtnzF+mjLRhyW8t091UUed0zgjqAqepCEB7EaI2QVfbXr0y+w5gd6NIJwlGAQ6ev+
WNInAgEPJcWeuLUx6rWEYiBkifdck+pM5Aqn3DQ4V7eHdMgeoKq3MAy5EAhZixSCNANp0t2XfLTn
Eh8dNlO4KGKCzVqv0loHpdyhguFwLiDuNmsf1V/symbhGtCU4Q1MDJl29ZK72JgCVNDzLitUwGwu
l90MlE/D3U+wcMyax0iQ2/hKFXWcCtTlq6yQhYgg2Unu3g5o1WfHmnLtA+24bsHuhSM2KmdhWhWd
w62B4aOSX+O30M8fJZ7wbb3cgY8q7KboRNutHCCiWPa2c845WSz+JZPoUdtsIUFZKAnpT0hXG6rV
0KqRgCXpuEApZl6fY7B61W5FzvJIA0XrbXbRWOpdcZCAXZ7J5MVXC3VqPV9Bs0zlPLnjNrpPZGVs
/HpolFTqMdxwUwnZzpTkkJuZ/vF0Zz5IQWdPqWsTyO2XT8b6Z91Ro2ZhlvGXsHb9MqTN5nu2Fezd
8TCXsFSYVzxHqQb2e8+GLQU/+gosd4n1Rh+ne3f9QZqqCLWOkGHbpuwB/s0TSXB8aXRDKqYfpedc
BDZq30mmFW7dz1NgFefduEUvUg+ymC1aEcNx6qrTTh0Yr2Oy7dWwdEUARDlDsWImBm5TJ/rl3QxF
abNi9gT+S4MeZhxukCEx5U1xM5mKHdf5xqEi3MUFmiRTnbvr7UZOtbM+CmiEvaTiaob63PRuknNB
RonkchYW9Vc7u4vMM+8RgJm7NUsmqTBZJcwoznPqdpaPy2AQbh281VuZxd8NEoB1r1jdA05KmoYf
4NGjKr6eqbb28ZaNYhLy5x4y7yGkLrASnrBx59IwHW6wcDlcMK8wNTNhJoAB09Da+LJcxdHX/IgK
2SuYqwRf10rA+B2HOdZMH8BSP7XiKx7G05YaQ39PcXF6V6tcXmqeYh7qTd656C1oyjaNheJbPJzf
vbGjzDi3qOUmH1LK/cmYZ4Qvc5jjFBWxBSCEgMuoldfJeKfOYu2akA7fJ6JE6MkjvoXjzoD+AVME
TT9+u4ldUdcrTJHn+Sen5ZkbKfpqK+jDq8Jv8KVLJKlChoW8+x4zionrjxi/eUtTJuBfJCMmFNHo
moYfUvdRCwZOExD1kh4UaNqi1H3PTBGH/V2O3mc1xuMHPqDZeeSh8qU8tPKXHjBY3BrQVxCrTrUS
+rizFvNxr5phZuTxOFpNQazJ+j65jVEnxbeQmKn8pi/wTaGoJzL82qUc5WW9cEsMgc5OkXX0Wpty
7GBfNZ5X0lT5yREMjQt3NyF6woAx21pEIfEgrmcBElo8B3bBtAROYFkqh5as/xHZaB++4tTgkDMO
+u8ktU4fJXGdVUjEvKtE7HrJ2q7/y0ka4UrPQjaui46Oo0azCzJWzDZisnond03+gCz7ZvGDAvJP
buBrMi2TIVY7qOznSnmjeXL9Jw0pAYU1Ox0vOlTseAfGKIlcwFbOEkspdn/6ugNi9lHNRMocMLi+
CoD4+SE3a6WtgmE9t3Ve1G3mcUXeh8/j3de7ET08nJMlT+fKT3ELhFx6h31kGBX7wX12pv2yR2TK
AKFZnjMNC0+yLLURQD90DsoWL6Q8TwkTJwaKs1hSgls2iO53lyqrgjywqArmQ4SQpz9ZBoKM7LU7
VwxG9MpdY3j8hcRE7GzqBSPR7Uczep1LIdi7MzMju3XWfWfgWqfwovlr0Og6eU+qPiIJBY5+uqAL
A3sG0nlQw5f9SWf8koa8TDZVljBg4aIT+Dd8YQPwS1cZG8740WQ9OMZ78X3NNhw9cOsaRKL4ome3
qXQaOb42qp/MiZl5KqTc+5j50XkL95nI0zQqwNuUYMWwGp+KH3wRHmbev+dMUfzqAGxoin3ptNeL
AwUbHd4UFYDataKjnZ6rmNSejHjoTSuB5cc0l4LmDVvsx5Npt4eqEEakJElAA+i3IPiFPYImrBhZ
a+mxu3y2Wn/dGvqYUq4pq6htjxpuemR+lIS3XPyAoZHzvNQW6i8kT4RwwFdmzUquygyKgfIFRfo4
dfmh3o/ttgrX/t9RGb0i/5rwbxhQcT1UyJk7/RfefCUlOUvHnZqWxQdmnXPTGCedT02BYF8dMv98
4Z5rUlYZIcszcbv3TKbdWRy+QTXJGnMLnTKKNUErMS86scXG4QSyTmNTzw/Oz9I5/rSd0bvoEYYG
5H3JzTc2Dck2ACOWbFgfH2LVFSFjj4BsD1YTMQft16X+yUwGV1V2GTFhtRZMp0k2vJ5w/awRa2VZ
bTE5/AnpWjWQ+sUPEh1hLYdbgVFdVjgPUOEJ5FvI/FbOcfqCuz7OtcPX49K9ZlUImotbQgPeJR9N
eY7woWCb/jnCU1i9T2PgiTDkCkZysLGElDCUeL4K6T1JGMNtrAjOqZscfz8PWuIQ5TdwNtS+aMg3
SpN85k66gjAUpqm6AjAYSAQdVjpDX0QRPO0QbvqAEGLlnP+e2xI4DayS8HRcKsnC9ppKMjD2HBHJ
v4WqqofriDAOEc6okjd2f7Ls7jxdwh7VQSXaUr3vkfcSc8e0D/pUTmg0zWVfNY1ngwskPJrQsqgB
5AJtLA32oYh3y/SONo9H9Mda4pfJhuQjTy8F47B420jlkHXUrhQa5Lemyu0nFApJ14kJZnhnq3iY
z/kZ/I2wwKD3ow/KjylHnGv3cofsE/968dPI2W/TEY6Lv4dzgMr09eRJRUQNfGjz+LHR4XEKYbm7
TC1NYWthb526j96iwU79SjBUN7eGiZgywxoLpdJNL/DnriSU8Hb6ZxFH75G9I/h27q69fl37yM6y
S6x5kZhn+v04o/8HWMPzg9ADJHKG0JaUoRyGmh0iB1Wi0w/Cz82ipMdkDVwRrv4n5IgrYI1dH8PY
8yYy083a2p71jGLXaXCzQmgdDoHcWR/C5sAnT86Mx9cSwyI/CSsfLxC11Xn7sbW7aPMaBRszXh0j
HMKTrjjEyiusNKWCnGcuTquiM19ZH8JyR2u2UPT8JVDWWvJcB98EPYLnaSnXnRIuBP6za4A1cVwE
8BXryru3zxEg24om1GJpnDDQUOwWI1/ZNUgdhXudfyYkHS5xPL+zQd1fyFq4wiR3K/wq8vDwfsQU
4MkxkcCAtEHy9KHtnuiIySWtdzuR8ILAOvhwCm+W/v1uMRwSIaDstG7olm/Rq/2IQpXV7TXzpTSi
31QCQi+tVk8Cz/qzpBOg903tTKDvrzC8eq9GcsZOlLnNFFglkhNKRh/x8Zl83A619nmgvE9RAWse
qAnLWSN8sVMAaD9n+WuyL5OA4TKPsxjgK1Wbcd1sD4u1FzBvWs+4OYKf1Xx9Wd5lEZp/msiQz/eG
mX8TXIvGQOdTCbve4a1Gk1eIQC7e33x9glEBdb6nV0b2hzz4QnlR8efriMnjsQt+yf/6CRmIXAnM
cmuJGjR1Atw28OWtWurAnEvxm3pAFstaxclT4VhyYK+FCYMew1zYm1beA9Cdm/M+Qwy5qjiTsWU9
vgZbL1fXYhM4DUYz0qb0rOCWeJq+hF7da12rH2pSd1jN9n2qz/AAiVZ8eVK//5deYv3BbzDWVJ3F
VoaoQiPlbp8almrtEekZgpH75Xew9ot8an8zRTLQ/5b+skH1QhQhSYS6Nhutux8LJctBJS+LxacN
WqcKNx5UZys0bhfZZR4PkiyDyTcl/lYc3y5udp0gfMx8PRmz6Oen3OoPeTZF1tjbU2hC3PawTkET
aYSXHFYOHNBqQ2jXU1cL4yxjccC5nmUazHHNb3ja/7gOZzO98np1caXx1zKmeZ1NEopcERbj8OVe
lHVEs26LljVFnZlxX5Pcz6eFPAPAVT9Wb+CGwyOhy0KoM5QA3rdZqBLnEudDGdDiZFQERkv6JOfK
sfMz1s4D91qBR3RG4kL55bWwKiGlVytDrZXjSt3rViMQpIMe9Ni6dbexH009fDesv2H6rC2wKXz8
NqMFHKie1LVRkz16gYs8AI3jE6DztvkmqNb0+2WHoqg95ZHum9AxL5tMrtl1vt5K/XzS9DvLDdsz
CrL13DbzO2bnelQF1HpFRwLtNNC6PDv+CK0scL5+sCMZPQwSgk7u9MoSNdEuWvePRly05WzBaDnJ
S6NLajWRNvXGkBp+syo2aSPNnuL4biyy+PSVDVUiQ38kiUHjZCwH+u0U6MR8busVty7m4nwXXrPu
XmpRiiMnSLFnsvaiTVkG0+zAQkGDoXy5RYh7L4trNLIhnIB2zwKIAdB6EbaqrBl60oWKKborRgh8
FGqpvrF7TsNl2XPjQhCjkC8b95UA3mkJgZPkiWYl+v2x3AyG6UfSDBOXCQgp2N8Tis17eAd6DbtN
n1OLGINeeP7p/XT4SvvWW8jIrfPOSS124SegPgkCECBInnxdLf4VOLqlZq9UEQv+4Busk6jm/OsW
XDcy31bFDB0OpUC5eUqVh8oO/rD3479buYTl6fPKINqbnOb7c18hDheWHENA+LjPjt3ibUCmIM0/
3LhhenTGFQXTqxT2G2adT50IHGZpLtGNUh0mhJHNTowNC6AWTa/opcfnT7kEfktBq5CWmBmONvE6
4eq6YUeASed/K+VhEahzj1ewAOdpJcEMcSe7C4JhSE0fwumTZWxouiwE0SQtVDaUr8kBlVAHYlkv
yYQtbLHdnDSieUcWzHKjCZyRRXx+a+F7kKIQNJZso/lDmdl1BhIBmB8qkKIfrSk4In+ZVHs63Dk4
DZIj7irsK6/EiYA+bDakIzAuLJoZhfFCaNrnNqLaEc0DbAxdOY87quGjoYFqZPXlepJ1aTCn4Alo
mKnfw1mkqa53AWV0wtxeHCy4ID/s/IA2mZQOVhhmaohMhJdbYuzsbC992sy2r4RQAOfRPXl+nfcz
GwXYiqGFwHMfJDtb7NaYREoICNEaT+6rKdgPfi2F1lQIcB/w4+FM59cmtn417rJ/mfD+mSbmkycU
BKewrsggJ7DoQEXvKyYVdUKdBbZuZiwGA7HyRFJZAtzhM64SRXmb6Xi5qbptz62OgRs35cpUsF66
abWg4GgzvJRFr6E7xAZCPCnltzSjJ3kEnADBqyZiokvZKcZ5qxxCd2mlIQ8CbQBJiujD7euS5JkB
zovF+BOMaUf5/7CNJhYyaoibh9YkCrE0KWEBZ6TpOb4veMgtB0495Q2hPQQFbRFQpfSlZBe10J8B
h2Zdx+RAZm05fwqxQiVaMJL+wSCRhSQ0WwQkE08c6AbDoG+hyg65/iuM3fayBtIjxcJ/Rv0NT4S+
VCnPK8s9yBm3ZDrN0eMJw6g7fk6VmMnOI4AsC1eIqErzU71jYpA4TDcU+At29fc0baVzhuQpxKGJ
bJCzs8eKP6vvTNQZ5V5WEXx0V+4IGK8cIj5GiXtd38nu/GwDUGkeOz5m/YUPCBgNBieGE8XGL2Yd
SNYdtOSBwKXEpbHbectlhWsdbt17tm23DwjpLUF2wK/LB5LWlwfS3LbR+JC4pG4l9ZLgk8AzGDz1
fZcZg8B1UQjNvBUNqxSdJwv0c3rkR1ZM7zZiSmZTMFM0G4BV1TdySGQqB9q5IPNfgAtKiDtKoMQN
HDrprrFPfA7kPjcgp7xO4yUnNJQ0f6NgO8TRS2TUeXOByhKSreAgdJn49oVoNGupPh2lNMrTxyLs
bOI9wteFLWS7YTxNm3Qqt2HJVoCXMlpdAqlcNwOX3DrfE1kNu8QXrzOZ7MJhN+i72NPpsA8WcN3F
zD1ZTm1cVr2IcNFVmOv65OgY5huTX1AdXUY9TW6wVydNZXkEot7eqhYMbCeuCkJR6pF4bDxNe2sw
/m/yZQwKyQSwT6pwa2V1SRs4MBU73o8F9ybEnieqLE9qQOuxSzFBp6IhJd3984fgWN09pz9ceAQn
M3GSCjLd2iI9c+D5k+Mdftzp5/TiCRA2d/LLf44c4dn60Y2EYu0wlFKpk/IpFMNZpYcrGQsILlQS
1fXlePa7MsPo9+ypJLCkzbYFe0OLIBRHOLOWaw2A2+mjHCsV0bczR1K47sg1ZPT7iNRYgrr2cnjA
iLudBSsBg3mx5ardF0aVaT9mIR7oQ0ph8WSylYmJOTKRNgqBb7o6R2kT5IxL38le66jTi6WgC17Z
YAQHP5LFmzNsW4MdKMTBQ2TENKmREYf96hgyCzGILXopGAWjTvTB/HvEsmGCByrNqdYT9Xi8dtRd
ilan2nMM0MzdyheziOnqvLWRDepPN9ILoEA1lvRlWcb57oTRuDx8GhFg6o/yDxBerzcq5P0mONJM
WuwQwjHPS6QVBVGsKQaPsUOxw0Kr47a56M1cAFa2JZEGRmCWI7YDU6rN4/diNl5MmmQo8uiTda3i
TQC7XBNqk1IFjuxXkEXkPVsUBQi0GrJiP91H+ysGB+2MR5a9a767SBwaLcTna1V1iPngj2vLVP79
5fzCaJJe9xsFvxZpMLLgsm9OYyLWNWKwy/Yfi/QNJmROrPoEnYCCL7FWGKPhRREdkBUGSFgmt5wi
8Eky9nJjbxR/Z2Yza3fmNB88C81PYHW4I8C9Ubool4+eZFpBYD8fdt8SRVSX72frpXj9GCWEk1sm
UkgIa3VCE88tOOaNuPOaffOBbFhpLkB6Gofb3xgsvbA0q4eBIUD8cu+FTvn+R9/3LUKVvXTZAPHu
bVuYMgyhogSoX9G5iC/1z8lolYchzrmRMNkwVojQdeMC9uALgFQVNYnqIrZ8X8xTIFeCBju8neuk
AwFR4v/PkePWfR8yZhgs3/MxiLizANahn2AMd3FnSb4Le5haz0zOLChlf8IqR2GA8y3w4trT8B7E
hHBjJGMqJOKduu5AnYivA71L/foMRaxgXp9KCb3CgypeMPOxqmi+9qrlAp7ZzUPFkGfAbzOA7omy
Kb1YtZNDRhpcnRDYMGL8m0XGBC+gEn1uORVS4PenSulymruFKfXwZJjlxEMjsDq+x6HkXB1myUoa
/ot4qFwaXkmMGDPfwXv1qD6HNRGLUdGqwCQdUg5IuTC0IFgJuxY4tN0RbBUSZ+LB4CmS11CiEIgS
b15zrPX24IRT8Hi+QQM68KoB7TwnsmWPzbCIvD/FfEVBrIe3FpMV0zw/ST2vK1O5S72YHbL7DlBL
3LXXAk2pr7LY3RQ3MgqaDVyrvEV2xOM6KmgrL71w8WJnUEMSUhk2n0tbvIQFuLdA4yXeRsUkfnhj
jxsTw9pQPpUAAsdwzWYz4xJCVAXnGnRdpgvdkl6Q38dlVmeIrnDN+MyrhPsdsLEsXviBsWoq79X2
UTQME2Rwz/nrczAJ5usJHveUeEDiZwW3J94XrtXGQlKa0HpEuWsyGceTzSu5jvEKNUP/pOju+/Jb
ZBrjunsoncCP47nJO5IPN7ypfE2XfvP8Ppg97lXyROLH+Hmk18fEPVqn9qaGWcZ8PtbJET12qPbE
SRxeA1PB+MTTzz+EwuQG6fAFe3ERGstLWa7YbJLOnd/TmcUi6XEuKfuqEVSrYwNRQoi/TR2BKvfX
Da88Ck4N2K2a7dDuzr4pxAEv8rZrZC3IgNZi7UXhSjV82KaE7IXc5V6t1bkWk+USSYbFxUI4C9XC
jgfBMTJgUTp0Fdvviq/LZJ7BdZYaF8IxlUZhtBeVl19QZXnua1BSXNpPbImCWic2Llq6KomwS9nO
nqyom7Jub/Trxzy+a3BRC5S0XwfW0p2gD//htqVAHQN48HWx1gycxaVrk5law/rQshkCQ+ruOZmt
LxCp1WcciAHRz7o104bZTTllwIYhXXZXW6lxsyIA3IlCM7vF9l4vxUDVEYAUhCgf6+IxnSbgbMhi
GfhSuKKkDxLgUTqhubhsGnYlPu95AjxMOyCcFA54PwZV3Us7i7fftPmzi8bSO69VSEBWzZ2snMR8
UI/IDHmuQBJ0ZQ0ZS6E6eeUp6OCPr4iDcHRdEthPA8UI94Iw9IQ5IfCOgn4pq69wdQ2gi77Bjy8R
gvTpJVZ7976SbC6wLQaMfRs6BAi4iraoMCSLa8Y5EFpi+/hjQ6HIZhHwV/O4K3Ns5U3uuXxrkFz/
4muX5VUSm81DZ7QT31WT/UBrOX/LJ7AjplEqvfUXsORYdT/ik8VczEh/R6ydVlZOFwVv00Z8Af+t
Uspaucicpee0RUcB+chu1ytD/65YQRj+CbEQ8JnT8HfGRPteEkQw/O3nSsdZB9xJD8FCADdtB1b5
gcFn/VtIunbCS5t0kwBP+JTc+BnF9iD9YZJ+PKZuED2PNzTIcvadTz/2JkANxwABwjD+N7WH93MF
kKSOnlyzDdw0NzHGadeU7xm3CFT+VaODAah44KdBXOUv4Lj0OLVuRQpHgdoKs5cVrNUurxhRa6ht
kcyreurrk+J/Vu5T91WvjOOLxjUxzJBuVmsZTmGfZ3dfOeyQA55a0UR3sqr6I6GLxE1LOz4pqe+P
espvorttXch4JXLeha6SU/mmYO/IRIlzejQVGzrLb5xscKm7XCBA7UZk23XjeHeKooiONxYX5lAL
vt5GLVaZ/Lx2MFnJaC8vQGw8bB+ePOz5vGkPKRHAm8e2rAwE/WuzglB2rOmMQTUED82E40CGQd8e
0BiLWRpMgUFYP4fsGDUQMz+uyE0rFZ7Gq7pTUg7lcghyeqGdqSWKvjt1/NcGsQAWqTG6YVfrMVoW
Q9smsoM9vYp/dUvGM+A5G8ElaRA4qFvQuMjuN/Wc/oPpHcVi4i9gmq9FSvzZFqyEYCTNQFsMrMCt
C+QFrdvB4H2MLYMz9F3pZ1RLT0K5M/fj/ZF/vbJON+xGkWt8LISwUE9DpD1uqB5lsU7p7nb4Pgrt
JIyaA3iLLqDgj1rcJcD5vSfLbm85tEjhj2iynzyRfQranwkxLjNKxpNa+6E6Q7pMYzOS/yK4rtCW
DT2G16CEu51S+vdqqeT5+TGbNhADToE2kl4ppzxYAtHS8sCShsj1AcwPi3MsN73/dHGEBx60Xjma
KaYwy656JHv/8IHiamD1kRl6Xxl43D9l+bv0O2HxUmh69h/sO4qpFWeHBVZORtsBX9Dhdn7wzE8u
m6ELw4WWOP1OKHnWQrPjrXbuYsXEvEQGmURhK9zXOkjRvOWUyVJwsL39e1QTXSRoEOJ22Nn5TdDW
r7NJQytYoRangeA+D2JwIDS3WvqJIbA6d4DEAbyqgNXSAeIr7xB3GQDdfmU9qI+ZWsUTTEFlpquZ
0oHzRUneylxTtKyKwA65r/a+su8I60CNqIcqFiw9bm9DQPjGiackR2i+iv+FXUlEOzfzJrEEdrPV
9JHSGN83XEuBPuzHBYSIxFulbSTniNvWB4Ho9jiA23k42i9YBIM4CJp2tZhRIzPOy4RawxCOs+tP
Zcr5DdKXoCFhCD+kL3VTWYwAgquHop5I4QUdvxuw+45NOuNTZUirH3pIFwkcXGgcxaocLe/iR9nn
FVGzWi1Ms6NOitQeg5yWisxp0kJpW9TCFTrVoCIaO7FQoGeyy1tlp1T89cj0roDAFaZIphKF9dSC
mHXE4VCh2xlok9vJIam9nNF8HEYZDvtggM+m3NDpDiqnEbxCcj2lGeYpIT+E6ExkGa5FilllCj68
TFneeWulwGeAWIKp4Z+p/ul2Y5Fcc3NIr5S4emzFLlhB+FAsxRjIu1EMa6T6HiUmGKK3su0CeSao
rhmjD8YrQbLClblh4cVLhJzmsZ/RhfEbR1/bJr+z2kz4cIqv3FkGuKDNotj56EefSss5/ya++jp8
DpVQFIReIWKhsD/YNh+s4oAzrU+e9FyEsBFe4YkeDWzfSh4Iss7F5E3B7jbvlfKcu/7i5MwN4Icw
Zbw3kYPh0P+9vedd0s8KQubc/eDSFBpdzTLHaednNHu/3sH+zI6Xi7qldfqhzC0iQmUwSTpzTi4w
Wyi2VQFBS8aG8V0dECm77+UevigVykIeFtvIhgM+UYz2QpG6vaoGLsqDftR1YAPQUarMSKsj4SW0
5ZfNhHoHZc8zmoejJzK1wnzkzTPlYnCrD4tXXkdQvAE5qUc4hqn2JQL/94g9tu7G9CL5pdm+DVHR
3iuj0qmig5wS4abHIyQsyaKZRDQ0MiUi8FY8aYU704p0qEN8jfiyGn5KyqCtapUlPWGHe0g8wsYo
0TYWpD2HE2iKHwUbRekHwrnXrQYIctfARybYAXZtV7frQDzFnmUfnRj2zwwXLYZKmNIjN8QSgQmL
CHW3UJ9H/cdCMufiDtNuntiBm69hNJlk87c+UPB8dxmdgTRZT0cNnvmi6ul8NFA7YLfZ1zGufw2k
7hU0xmgSSQFljmdCt4H68LltqPWibhDrQ2fhMCrzt5QH2QAFkB3T+u8WfsAabAvY+ckr7wJ/PnoK
MV5cJiLjVSq9k7YXnVcjhxPNOQHuotvFyXd/Kfg6SrG1wIW3eG5jUdgsWPwP8cjgeWQI5OKUpYxA
38ZapK3Vzc5LoTSXvCbuaNYS/E1vVe9g/qkGF6mgs7LsWbUOWkeYMSYSJB/bO+Yxx70a7kjQAnQ7
hT+qzwlapAFmBhM943mKrZGDHxpnDpr5jM6Bz8ug5dqfC5pqsVRKdkYUhXowCpsoTN3pp3jI9pwh
bjLzOj0Xs/cJdJOvjL8NeaH9Dm6hm57Gedm/8hT/1gGMsncn0wmNeBdCHAg4JKmq2fO1b6wZiTnv
E/oP8cuJyFJ2EnrPovBk+k8wNX8QoPmL3/ybNaGA14VRsVLrgXqCIFowSM5TQLDkl+PG8gUouSUy
EANbGwi+dmfdHaMlICOYnsPB8R+T8Y5IEV3KV1gLhX3/Ov5gv9IgB3G1ylB1FUkXsitdM3QGIui+
0EGCL3P3h/TBoCAOidLGq0NZvb+EG7yCflu6i2C4GBCRdi6C8NuXwmqQLelv3GS9EMlov6TqK2Gh
xZ1t+f1etsHXkNHZX3K+n2LbFmWbaixzUk2I1Lu4zPlbwek4imaxl2l3DBcWwwP7uJ9qQzhbtkw5
OQOr0+0bOz/CjEYhUZNz3Ukec2EYsFq3/BkO2Nju2oobA2q5l81d/3UaolbC0F7g6OsIKSta52+H
ddTkUIO6eYq5VN3us9C4Xt/LxubxSyMGuZfSMkq6e2LzTCDAix6jxk5VIsFLdZ0haD+UN+//0K3r
+ZPDjcLKCxda51o8mYFKsQ6HcKlGoSN3zOvDYb2zri43es6INHiZnqrJJGkk3+c8v1Krtycc9pRs
c7E1cYsSX1tnQ47/rYmjEiU8FjFGgUJqMu7qgV7BpmHJ9Yd9gO9jcesnDUXluS68bkKj1bDuc7vT
iEnmdnYkCwG+R1jkROI9rBZCaS4cZc+LJ+5t2gYTq5xw1cqO+1IYUtpIIjn0YtXLLagpXm2nhVqs
d1w+1845uQlCZBxma94h0LcIuLwcwCXePIiU6G2qjIUU6MvryqUM39uJfw7inMFPPHYMU9gmFAhX
jGzg/WNJeAASnD2kxdlJGvYgyYCQJoirc5+skzjyBjk9UY6m/DKFJQHUpc0npksQjloEgT0y938L
kGRQzwlMcQcSSNgnaYP4efLQoLAVpNCGH9/9XxdKHv/UfqlRPKDLCJHRvW8cWxvLFQsfX8BZ7Uk0
BMTTYahcGOkFKFz8dtyRPf//1iszMlbwwiPtHtlqCbxSSp26KthXIP/HuDu12OEF3Sv4PH6h6skv
jIrKL+fB+Dfxg5CjAy6XFRM0WZdoUiQmsa4Y3u7IksihVWWGKQQH4fhjui+1ypPLyuWYQvN4QUEk
vVmemmpOfMwVhoGQIzrWhSmGxdcF9M94o/TurWsCJOOCqsHfY4c7u6X0ndWGRLUYYZLQdheiF+Ir
pdCrHw+d/iykacaD7bjLmrcKwhqa7EuQF7CbYTfVZrUvwEWthaHBOw0U861GYYYonf836b4esivX
b3xvLMYlnrezq62uHZPlJGuaJVd2aFPPWk0xOzmc3GGjOhA3DUc9xK8CIX+a6+n7fh/FL/XNEAj0
5zS9pnrpNrGJCPZtwgyUtuKDRAID+SzOqT9iMVMtzyZoaqix1+KfKGytkHtTSrTMzv7cc6pfEA3n
h6oJgKYXIke8bp2yq4U84Xzknqrkn06yVVF2W/rl5hM4yCPrFqYfCvyP2NjznO8In+5sJBT235sk
HMoQIFnadgx9i/jyyhgwle97qoeza/Oe7r/FVgnJ6MM/BEd3+XUjqFaxL3ikPnsErxuFf3hCGMWz
7KaKe3bA2WRTWVUxtv8NxvgmTNTcB715Yv2ddDr8sX7/ojmhj61inEVRGVNs374NpToOCYsF1ZIe
KL4ZfIEUkyAL+yY3FH9bYdwJEM7achfwCzj65SG5eAS+nI62MP3ryzpil9i+6z/a6Cb5SYSlrPXX
NVrdQNz5uOZTDDQVMsl8rYKx8kYXM5+Ys6wWgdnT/1ADad/l3x66wvcOW/AuGQhNgM6hICUfcHy3
AetNSTWKZvDILdvJVFmOjfFuXnacOySgO3vPUchkHIEbITy03oJW7lMyGR1G+2yE9lmj8CTKO6wR
PzCJy5Q5WWuiV6izKWXN2zRumgAuRjQCDGuU44eDWd2ddlM3nDMddd3mNBqLsDElKmvoNWMQ2mBb
nEHCPkCKRmTBzoe0Wt5R4CQaUjlzdOeYwCQ3CnxPeg+zygEM+peDrGXRQE2JitL/4DvU3NIH+QmT
fa59vefXLJ+PAOK6TyHoK6TfwFjZfEhL3zBinJm80Y2n3DmC2NMojcLt+9B51IKbE1XLFsxYeScM
rPI9njEtUg3IMw2aNPpFEwvnT1EBG966Y6RG3/FFsw0Hw/3il9bC+Hsrj3Z+9T50NYMJoKXFReeW
4GEM8KKNrG6NM9xvQbuEtk49pPW5ggDTfB8aW8zR/Mm2yV3BthWe7fahpGD52eoWI154w26LZ2sk
tWvJLIlsPRGQU4/8uBYHDHLxiuHHvzWrJFCBGs8eyvxoeo/DZyKRbtiOhkyIuK45j9EbK8KL/uUB
ef2i9sUxNBo29X4zVg+BBwl416IY1QE3TvLz/t3cJAB1ig7VfRkWl1yGnMMJ1Lo30KE8DsEyPIg0
A7bEKT1/dkX2U5Tw/eOZz1D3Po4CkpXIZzMRWSb4qiZEVlMkF7jUbRIqUGY09yePt0E1pX4pMOUj
d+akBcBLP4paMc8Rwi3q8+geRmU9rj803kh1riazUqszdOOyiKEoqX655HeNDyhquJd5vR5QYHeF
FOi6EbMoi/rQEycvAH96FII87JIR7J/iT/ntPaSBSu2FdBLBRkS8VMNiwnmoY7NhKMbkl5nUt/3B
UgrAzRPLCymgI5vtmMBmmhfey7pMmZ4nVtlF2d6V3GRp3Go3ZiOy277BJ2WXV6YW5C/7FWd/RZy9
TYPMidoePj1KSRlLYjF3l6AB/PtivjPBgjC5trPqEmfqIrrbWT7+Uiqpvlq7rpP80DqA+44RvYZ+
AdFv+fmNt4jjnBkYj06JSQxZkSsZV7YrvSDPK8p5FfJVi7NlCba7q74ToXqrvesLymMTYt4YxBk4
WLYLhrxLwBjj6KHPEnEc2rF5SEi1dTBIb6/bkp9ZxH9dmAUaJ4Ny5fpcdT+/X2xfYmwlC4xwFGnA
k74t4vqzUsCxXfvf8RWRBoo2XFNoTJ5X6DiqrJo2NfejwysDLsv8Zam4ukuT/owwwXbgC3P3vNFJ
A8wLo4QUpjdlWQI57EyrC9Yh7iMsxc/+Nh6+2zSsvw0bHByqOYIpr57XqSunCFYUdYHpnaUnwDeR
ZIM1VoqZYt455IBdkYt7o7qu+2YuU5U+2HPxptfcFPJeomScI88XE8h+dTcvH7Sh5LnzWegReNs9
IM/j+N4ehIErM4ZIillkhb6y760agm7PD2dn/pUkaT3avAGhO7f5BWgqCTZySQQKx9OONRgXTyhf
/5RIaJf1c8USg2y8xCOw2ji43yi+DU+uE1mpvzyh8STO5rsWy6HAy7+J/yb7GpdVqn9JGimzVWab
wUaOadToqX5ks39FB0Se88h/vfGo2CR4PdmuCCCd6sQh8yFasKXFoR9aWGVTgeN4fBqIM4JKFMw9
t3qdzqwtHA+8dNgQG8w+XJNhs+Yj6vj+F38SONX65fww1c+Bu/0yRq+KJSWzhvSbGITHL1wLbH6L
B9mQLTi7DvwrCA0ww2OrkJqOB6oTclenCOFvi2u4Oflm5LOjM2Go9GtUc0cvbtZLmFu7NZqiN3Fg
N6mJlzQlLdkrHLdk9HX/pgIITU/rURTwlfhZZn0dlxuQ+4wN/DoBNQM7n2DcrjmYDqLljKfYtKaI
gkeI1qsdmrMdSpJ0nOd7XZn6xlE6KpH9/Qe+8rahnMfYnJrbPQrqY1gr9ciuC+1zAliT8qcGG1oh
RpcRlaxA5Z26ZJEdVM0oGbXeVU0BO75i8WtYTy5Bm1R5wf+vsGEVkyM+me3/5EIusiokRGqymSOK
2S+uNsY6pRWxtPCmikLRHfX4BgXbTf2EFh6VTt4H/ek6LXLIyBggaNhYkceklIYCm9mb6YBmo8ZZ
yj8fWtGvdZ8Mthima1ifbmmDC/d6CKzhr7+P5jsDfF54qoSWi97Bwh3hvoSxULtQiYxarY3QkKnx
zUINZtUsIAXCNVHzrY1+AgCXLAgt4JPTZRzqIqvVuyYvBxLx3mPtosUT6rIGRcuaGX4hXXqzC4A2
tk1YwdHVCxxbiSyetnGoPUUAGZJw116YG+1ROv0K4ew69xjMuCyDN3kHV4lbG6foGSCC+/rjlcRf
4DRivLx6Y9zPUEbOG/03lcc1CpM2DnBU/dcsdvDGzv2Xc7VK9dJ/8whedk1YfGhM2dim3n7voUw/
QwC1lItb1hx9qg96R63r2un6OK6Dyw5KW04PXy99avPYPAZBxsjgR0HUFrjnlksXeUjxFzAegD0z
yibwGzwmXlZTNnHEDe+2K2zDABWaCLjGfjkYzXMV7U6x/4vtXOEwmER7stctS+DNqfA3aml8SVC/
x7NLeNxZ6++HOx5GvW3C9k3EG0IYqilz1cnb1N5Yuu7qHJnRbmBCkiXWC7sqzzu48ZXcuMlIsn1I
kPRndc74Ndh1TWyKX8Q+n2PFRnyZCXkA98kvqEBzetMLzeepSP0+faY4TkPc5d2mAbhWLjAnYRS7
1s5dwUoziSn4jc65bAMJjsYS1EtVAFlPPOyPkYZqQadqXjRfOC6mgmIouQBNP64Pocnz/Itq5LH2
ggPNZ3+AizyEFBsf+UM+5Fz5GkUcqYm+1IEgQh9oxJWo8YAoSOIl7p/xOd1I7g1ZVEvDD9becBdQ
rKwzSiFvusHwlxtMDz4VTakt9ZXmqvOCl3IB4A3/YJmMVGNIijKfRqZT72B868rbfoHT0PwUFANz
7p1Kpty8YH3m/f0QPyEbA8LjL8vIMvuQqe6kw9N3L1XOgRyPk/wea7CwZfWCx2J/yzavYJG2rLST
MiBvhfZDydyAfyiaZQSdgnsM9AyUlfF3tXHKjVXu3ntIEeRWH1lLKVdwH0cVKywTxJLkIQegfF4e
HriM7wXzy/R3R+Waa1/KfeePr2/IPDnsJRLN36H5h/QT16CtVxTO6CbC05YIuJcprINrYIqb4sI5
uOEzFpw1+Ul4k/8MoE+I2eGLHmv3A3fqP+twh3hliQA9fI71TJ0R4ePA9esg8AfkqqeaGUWydXm8
0xaIDYpljcnBWSi3sGSU052pzuqEU2K+rZWwW30gFzNP7W8fJgCh0QQEkNHWePzN3QLAn0JWghDT
sTa0c6NWxRLwUyAWkSwS1x8iL0HcXQc+nBfgrWnrI+y0Hkq4GvBWyCUNagmRNl7rM22gFkPAtvyh
SowXUDR3U8ncYODvo/CwAEQOcOClXkTAplvhMbamicyhGqvzHO4pa81wEuzkwUpgFNx6Hc0QkyaI
yED9gxM9GB9eDemeKnoaQAdKYNjofO/ZMYDps12LLwyudx5d8Go4OWS5QZWYvV7XQ8jqMZmii105
sZPqkElr6BWHwzNrpg/BqGKTpElMh8DVYkV8XIN2u7Btjkb+eWi24upG4DYLqm/j2x4WSojnr+BA
lzwXmKn7drBbkkg+6GJ8K+Vt2o30gAf5/2D3RZY6jVD/Azs1sUpvJo4jEWTrOEhdhBmv80ZT5UnI
iPfCoVM0VMicOnPZr3k4T+49fgaKt9JGg+CxyQVndNkCu5DO+E8Wc48t31cgJDVWjpERaWjUAyxl
u/hwqzfl/fsCvt2wWnbdDfw8+WHJk3M1mJ4EppQ/gben/aNW60bVkFr2lwfloKnEHVkUUD3G/SeK
LF8Pi7LcE0ajQwDjNCfGozicHRruBQ9cn3GIEvStCbf4XUSNC5tsiS6XKbqWaYnznks1QBdpjLqe
P5RTcKT7Y9NfRxDnvpsKATTkp6pUO9ic/qmb08eSlr+HWCYWQ7m1/Akkn5CWKhwFLsa6+71jH3cZ
KOkJ3USkWvMnNq3PLSur1S6mLqcYhsk2+0oWUHhnb8wQyCk69jWo5qYIiVJyaPzsQSM9pm+YQ0ER
4JUVKlEZ2eNivSPO55X3roXKPKDWiGBkQ6PWQBKhyjpUOX4ZLq47xC+jjYlwmrfIjirLstknnVoh
q91UJ+Y/ucIsICkxyud/S/U1o8/Sscv5+R4Tj2cf3iQgkr5xAFW5qtDOex4MmqZ+1aI1Hdb9xf6U
QKwx/rHotWIgXu/Rkq/y43PokidqJJqyOHpvfJ9sI7LYIkcO+/Ch3UAcETjoyGL62xxSFrrbEVm8
H5Dk0y+WLTglba5fl6Fr5vzcFZpoiUuRr5+wV+mEV2NXn610sTBnEM2+LmQXUDscJk3yMK1QvUL2
GhSNEa2AEi3opAwHjuTxuGim+R1fbyFP93JEr9dUN4SywlEcdqBbDhIGh/aW/S7RDMI6Lax94J+Y
9jWOeZs4eWV/RnRxNzi7tXLI4tTMcsKUfJ0wewtXlLZ9TEpeRu5t1zOi8d0S0ZisgvdOcNddOKIP
hnA9C0db64H8ATNLxHT7aD4ykfVoONlNMGcyl2s3iebLKsZDbZx4PiIK8NcF1qgsk85c2hv1joxJ
iuEFuUTE+wN38Po89Hyv4lb2uL0n2/QXhH6coeOPDu40TYXdjmt2L4yOcvAD39/0G46ksnfdJvPa
YpDmA8BtiuH9lHB5aXT6l7ViUYpnad/PJg89fS9/Ev4RUbafGpjxxAoLOrkCIQo3R0FyZ04bHybT
nXTkfAtOj/PG0DrDtgdQ4RVbmqVj8F1YNPJVhvAaRmp9sK6tcoD3NH7fobhTjCtSjMYnpYp57WUm
BeTc5S4KHGwjjHUbfYsLlTfedSQSfKk0klTMnCKgBfUw9lWQSybAc4Hwb4Emfii0/msN2556Qbvk
nX13joooRNFkWpFsC4vqPFJ5uI2y6FGsbqTQHXKr7kAs+MxKRbWyZOOicEjjG7AN+x8SxW6fWXmq
EGwaCbBaTAB0KBItb2kNnVKSoeJERdE50qFMGLFCJvrDyRlXU2simhnlCwGp74t53yVA9LT4hNpi
9ZW38dU8W/PvnKGtIYa4Ee558bLovnfdjWo/f6s/BtHidQr01ikgmcS5ZHV9C0pKV/k4e2Aab2gJ
3vV8qzU57LCxLLgbR6Jvoq2vx/pLnHXaNDYRTbTXINTMJRZZkUMkdjI0m8llmQyHIh/xItm9AgnH
FQDc6/9+Fd9tCYbtrQhB2mRsirGP4VC8b10PECdHLREPp7gVx6qdL1r+kwGomoIE7ah7z2lC6LdC
FL5rrMFLuIHWMrVjYKFNThulQ6w764oD3Mk+cURz4R9xuWP7LnBf4HZGqTaUH14JksUEAKeqkt/h
52OOhvVOd4R09Y54Z+QifyHy52nMH/7OhW77/1BriAudTF+5vRwptguO9S4ZICcsK4SWNzLQv6C4
ydeeXwOoFGD4wzUK9alKdcMhgSImExuaxOPuLB0IGgbX5/cX4klfjsV9/A/K7XYz3EcL48UND1VW
rW1Tr1ON6JOxi+DP5yMV2rp7IfFP/+dNlSPJobAtPmNXM1qfMcHJMvjnygn3Z6ztQ11g+cUk4J/q
pvdGcGZidlNTLadstUqxGMg7rcSh/YE/fefAVlkXiaECt4nyTLOJpnuT3gamkjWtvhBSigCJiPYA
3rIIzYYtEtBaPwzUjo3HqFNz4+CxdHRLB+0ROzXlv4asnWbQo9rjiPvbKX5fZ8j0J1iSbsRBwxjA
ibxqOeKgrKe7Dlb2P6R6R6xAOZ8NR/ITYvTf7xTtt4k5/7fru4H9kQBdR+C2jtmC5Dcbdy4Dma4u
7mSNXPGtDkDyzT9Ozc6a2Hr0T7PC3o9R7elfSFEW3OlRySo2ls7UHZ+zvpNfIYTo6fIfojl/FN8v
weR/cCKakPCXkRPnu+aJ/actlrja6rS/G06BOowVeA9tg2i5D34pdZvuDq/hykq8eI5ztL2h5xUv
BCnmBqNIjYkX2w97D8nz/UJI0Sidw/sa9YqDRVPNyfUEJSRBXRfGtVYEnPyP3PPp/whZbGicLmYC
g5+LIFpdlxwsuXru47X4mG0fQQQSspZ5xs2H4zteqZCWG5ueftUpWNPBoq31OQJfNC9L65+/q4ZZ
YYCzqGRbgEgvQ5WJWLcM++to+dzT32Mmfr5qbhIPZ0n09IynE+UwojqKHhU9MoS6XhJmxDrAOFf+
Q7+5IGpl06+dNDSYPmH9luC33CLTTNlxi1ofJ6qiOg31Hw5IyEZKURtd6XgDpN8tqXi1C1B08bL8
zEcQaNbpZlBhkA9BjUcVa6qn2VaYItDqLJzTwKtXEdHmLBYj0Bt/CzV8WjnL/Dk5gBYICqCC8F5S
Oehs3Xu5CT002/2bYC0Oea31M0hHe68/1QjXdBSf1XZX/YjIdLQPdDIIC2kGoCta8bZKz8weEEn1
02+VwRPakOHTTlxh31vHS0CNumLSULgJ/ni0JFVteZo/Xi2nYMYNBPZm469mpUAmKgq712WgO3xq
88VKlwmSxbIKZRwGTUOvTQbhs2O5vtu8VBW6b6G566yu+PZTFFBZPozxH2i9t1IohXjtwIYts5xA
GZSR4TlnYi1XHtSrNIZl81DR8L0REIKd/xNKaLaLVEd0k/dcAGyKhiMg68Jpjr2AWsTWEpviyIEG
MVw8JE5EBzRreVNMLG7prtJYgHPuRV/rjoI0cKbEyAqi9MrNMXzwKtUVl2EgZ+mNmtXsquzmwplu
8RyKNNtSKGM6PG0WBGpzTEuwQMHS1GolKQ/Z1URSuUW0psCiJZAUy2E2jW/SQ5WjTh2BOpMvExFc
gvuh8NmgQkLUhIpZxvArib3gQ60AO/+QmKleENXXgl+jJ5Qwt9HXSzHqxqQhgveKKg2jAl/nnRH3
Wgq6EARw/CKzRZ6TbCK3YD1ilCJjb/6qilHCT/prBmRYuvp4o415ceS9YJzIZoIeqmEAJQT7MyEM
852JJWSHLcJO6VKSd2iCkBj3Mr2RVKrvDrUNaIC4ozQD8AvxKwt4bkq9WBhcoParh/qkEOC87wfT
XvEqu/7lFscLdj7wrq91tJOYK05BFTgSDXAuCB+iv7BQ6+j2ou1xnFgCwojSwzOqampm3QWFPlmc
nDlnGC/21wmM1Klc6m8mE0P3lLwFH2AVWr26rZYSNnAanS25Nln9NcUB5EKN21Oa1lX13Up5iPau
+9Y94GhaZP4kuNz07dStuUtq4fbiAv8YUFh2/N68IeryNNWsiarVXmRvXguwvy0SX3+9ZTM2/BTy
esH6ymu6TV4RMpoGsKRoCmq6cOCqj8dszvgTu53Y2wuYix0jZIjk50pjNSXxfioACjHGyBTkV6wE
DKRdhoanoO3DKVn47U08NZllsV0JKUbsfswRoqhL9H9XhwWxcJso2SbiqMXCWOZnpskk+WwgyUmC
QtmU/8UVfy0lrtLbQrVdq0LM60VEXwb4F8w+nnGF3LpDpXmAc8bUEXmw0cYiSut7xyIH9DI2kiYR
fzmsNO1k49pBzV1SQZJvg0Cr7wF6LSWw4RbaHTEwv61s8JrtUKIxOMa8/rhzK2NBZa4ESBF0AB99
Edcv0ev9YP4bWgT3CJidpuJizkcdwFr9TDBPgUwbbhjE7IKm9u9Np0RbfKb7hm0oVBLUmSxzt0wO
nlIwwKoc2uOCZG5dcn+teb6jQCYh6ebpmtZ6OFQSpeAQIQa7APE3fsQPRvAdd7+ngg70o232rU86
vOaH2Rv6BDMXLbyThzS1Cgyw2q6w/MvvRalcb5+NO6riSURN8SNUR/8trRuzhMPCBF2MR67mozFs
wIyPXFiiNhNovOCTjMvcWWaKEWtsZWt1Bgy+NVpBSvvTR2Hxoy1lT5vSuggmb43F9kSjtA2XJ2Dg
8AvyRjA2iwzufWMvJ7C2mw1YH+ljALo45NSiNCXh64eWP5TdS57zQzYSm2AtDtIuEQtvgJ066Tv8
B0WJwWKqksrci3qSUKTobshJ54A/YUdt0sJRB52RsITz5zvetxhOQYkUyBLUxbhJsObupjQnNR/m
1XNfz3LwPiv9Ho1akIN22AWFvK8r/A30bgnxlLnedZTMghmnw7T9msFmenCqvmgz1qXKw167LENQ
z78oUOBT84FBekMwn0ZztorwQ2p8jrDXCfdD2gxSbfbryEU+wM9bKlx8OHhXwWj//TW86sZ3QYaX
Tw1Hao6ixBpCbL3G6411639qRa8V/7ERXWJUi/OB9feTFMCpn5D/fXgfqZKkaAKZtmxoDClPPrKm
TjX46fKYqCL7eS+Z2c86/VtSxaZo/0v5PqTLIC4dhz91hBk/tToNqvxMqXMD5bROs3zBpPPtFV0e
92SaUINJRpwKQ9ryNkDuoqAdkaCi6rDEw1Vsc9pXbigAyORPu7OipmDn6VtVktLBiwppkje5DfOZ
NvsAb1y/q26iWVNngoA9IXDHFdyKJ1jHrkSvoDQZIjksltoYX9HCT4E6gWtUOlWgM/k63+baPJSE
+C7TFuWM8sHYfeZuqfCLlvifeV6sO0/nUGQlifr3iNNRNF79GFDi+B5Z0+5+Nk1jkZsZi8ES0Yb3
PEiF5sVSfWfpg0Cr70SsfOZE3DI8seE31zESSEJXDFeUxT86pNLzpW1gVProxcDdLhTBjqQT88BR
Kdx7nxWHLF2OfFfchLmqrXt019jMP7HUKTyLEK2f0vwLuOpVKdnoBkx/T5X4mOVxCl+U1yUA9M6m
ezVAabSBQXo3rEzQehD+ZwhXIIN19+RC7eedfJUTYmk0e883XT68jYZSusxn6FvvEGU91Tqabgm7
Pu8ncpsYdT5pH6NvKSQ6JmI6qm1f7f+hKS3nNTeBr23cisb4P7YGBZgdOXrCkKl79af6eOv+rZsj
QtE59C3xSibIq6Z6FALwYNlcz3UJNUg9HIQVaCXjmu/3wcW6PwhgcQz53HTrGmpyE0oSCqp7FldH
WAp7TVMLIB6p5aEKCkRIcTm5m5VfZ2aqj7Qg8TgxBxk5ipVrviHqmqx5o3hr0xHWmphh1ET6si/q
Uxu/YsJH7v7y1lB9dUSFKm1NpAhtDSnNT540AeteC9iv0yjpO0GS6V4XtbwcahoIt8pbDvs8OZP5
UhKU8Oe9BMV+EqXc2OE9KWF9Lyo7N00elSYZ4SMLVUST71sXA6czIO00IK90IH+ZLOtC3QTiO7lN
BX+t2CJpp0FbPGpAGbhhE9iMI1fuxD3pyI3+dngtxpkiGjIi12VKmDV1fYYuJVQMRztwRTZR8IHq
11CaMY5am24sGSswPAq6VjqVXxvj05TXp+j4hXhRZaLuvN9C3FuCZHQLAiy5ekTGGxLqq58DUy2r
Q8MgG9W/x3GUZCGEXO7aJ3d90hFjMFh7rrO3wPQ6Sa64EO+mvWt1twJ5SJZCHRJlgEV6Y068PXXA
gCgiKRIqcCiFjQf6Cv7fhgUbJP+PzC9JujKaTH7jDkGv2yC9s2wzCjusQO7wNOgren9Lu1qc7aBM
hQ3MG1eo0Wvh11/WpqvMwdbJFOJu/8v3Jw01VqMf5tVEFjgGnc9Thc7ArD3WEPoHHXwi9Xjptvin
hnVU14scGc9/3yURZ/aCSIi7ljmyv4E3Q8+86o8t0LIilNrW8L9uL//Ho0PhuYMS5Ni/ddCNUtXH
plEibEx/5a4+3hY8f0pPZBPbYVk0bqOm63Sym60hYVPVYDL3ywuEKrcTaMpOSS+t7jdBPAijYlhs
6yvYWZtEa6rA89sed3kOOxQ5lp+17dAodKL7JDc3rYa+u+kZj7Wk6LQrWpDbG+gvl0yakuJ36yoA
P7oKAdEmu0yEqd5SqTfsQ775n9Q8HmME1twyTPx5/hV87NqxKCXGAtv3PwYeCkcPFKIQihZCe4p3
d/NDui6UnW4FiewJOknYBiaAqdXRQUdlG4a1I9g7tUjOwq+2rticwy2kLpz3IsTMUO7LoT8OF47e
vS9ypaosx21wj3tXdyqX9AMIs3/ao+oueHQjEUhzW5RlpOPKjC889MS3r+XyKE7rvaWN42Dp19wx
k872bbcEFjIr97jQq7f86pvWvwf2TNWz+42SLx9h5fabdZTnvHNv6DIUpKYigLCKaUOiRzqCZiYL
0iG0xt8Y1nSJXUuJ+QbG/QXGbCnK5WqQWvd1lIPvS7KLmhA/fk0SZh8AFh1lTIVF8s0uMYAmSFHl
IzO/5M0GrbDjqkGeuSAH/agzNx9vD/oNrcEDX23kSbjlE4aBXkqotpXFqXNi8WooAtUIEaC864E9
/EJ3ki0VAUm20QBu6Y/2aRZRmZRkkQwjPcvhN3uEVBIKLkhq/Mb/v22lxPXApSCqwpmdQiMkXi3t
+tbd8YTNFjuGasKhl/mXQpKofL61VQ/5Elj+EvUD6kqN6wLdqP6eP7tBSO7KGFJbIOMYBu/ZTJyp
3vk3UJXNTk//KMPWMuMjghgy+k/5gQrXosB7jnD28IXxaLku2dBmxeaJn4KWaXzt/k1dNIuqdstN
QJJNs4t8I38/XJiCFb2sCUrNr+AGuXBG/ul6BgijRGiS0eohIJ0uwBUJClquMqXX6WmroUeP6OPb
w+fg83dCSBaTnIx9n17DW8bO/uej/lE5NqXGIw5qnf777/8CtyG2dad6NKqu+W/h+gM3GTSTPPO/
1V09biY6yHF5ozyQsm/D8Vlu2V+9n0ccP1yzy7e9DhpvThC8qEkFzyJcaltEbJl+dY1KRlQu02sC
M3KwgK7N5KHNNo2FdDifdAWoR0fpZ0p3mYR1VB3cX0yK8X1yDixb55zrWqohxbAVA2gIWEhHLuDs
bnhB/puffRVKvbX2h6qZpwa5UgUdVrV9WoodAOm/ZgKwjdJfnyX3i0ncjW9BdxrLV6uCz6/z3SH0
W3IjfQy0AaMjIEx5QGzkIloLiD+IJ0hsNwX7P/2ZOVain8vAa3akA3SpEUu5FaPSEa5sfQ4O7ZlS
y/brNEUh1MahGYmKoMKGnJl+bF/3os/FvCcvfuc9uu1GEfyCq9hjFmTExzKWCmKsWI5mWPsKMVt4
dThewe9vQViCuMqI04WEgjqiW71VA6eS/0t3B7Gps+OLHDpfBdN29ZnJQp9BOLOpHRSizx7dQ7y/
MxDIC1Z7axxw/Ja6qRqy2QIHnEYYz4qx9j9JMwETclnMkuQW+qXGNrPY5EopAMxCZwab3L6pVef7
ArVtNmG3YOAATbkgm57/yIQWCtZipoaGuqYAQZ6F4l0B/qpoC5WCtWWH+KvtQQ5MpiukgN93SWm9
5xLLsr3bia15zhv4ABXiSNQfVQyNrq09Iq3YIE7aBTPCZKoZ73EvORz3vwn85M5sxbt3ZDojivTb
81q6O5HNiVc9ENj8sYov1xxzeABs5atCAy8NOR/h4RwdH19oVxWRxXM2z/n9txAgN1FUuzzN1pb2
37UTM89Pb/gP/8oMaPQsRjaswvlHW4U0KBWAlCt2GBhnUvPRfaaxHDVj58nmrlbZN4bGHdoVQOQI
x3OK1hlt2mukDhokGkumeMF6D5lsHJcn/jI7GvoTayR4fwfGLcU9iTMuMSNQuP7UxZpolsTn8lrl
PUwrRNFTVhflDvbA+ES0QBa7Nl4r3QoMd++uBDkr3h0HJ52IiqBZYUkbQIS2XZOKZiN4/KbaXnF9
sbGbab8BcHW2v0MSRAAtaJw7SmsDwmfSF+EbwxAqfooPJIwqHrsVd+/tEXUeLbO6VTCadFc1qq/t
rEl35w9XBOr/eGbeshoB3BFYHCdVz2klZVzAV8NXqfgqbzTcMjVYdwJ5habs3/gbIZHG9M/RDypp
YP2UG0BlVoPq0zhgPB1DI4QS5DYu6PACl3SkpB4Gi35wASL91sKEnWNY7+4+0OmPpr0INteMRvzg
HDzMIjCD/OWAknLg7aZxSJNNDLQuqdZsam7u6siO6HTX6FIutV7Cbxd6SG1ILcjI8E9+DH6PeRqA
ugog1BVq0bBYjCE7jo/eMCqInxsJMhLtJX5bC6fI1tOChUBSh2yP4puUum2vX7nId6qsUKWsoSCy
OxuoygkkU3PBa5NFcKuF5azm/pMMtgWt9s5xxtu5BIaPK1+1hB19um3xacIb32Tc3v6MV0/Nz2mD
ErRaFsH/EmhrKf6N2xwtuga5YPimYHqLS6cPGWnaZCebZES/K5MDYffnjgY0eq++wD1c3e9KRA1v
D0PzLgD6axqr1Zh+ZiaMTKj3z+6zldzr/ysJeP9XFYbP8NJmfLjAZFcbSa33swFghZkYp7LPy+sH
6nEGkB9yKM2XVVmr4D0HT8bNqlHPMTRXFryv0wv4LkqACyygcXl5FvqP8DH+drGiYqnQDcgUD1+O
Mb6wuvqoJAV09jvGOkv5vydP1memINmt0jnjFkleKcAKm/pf3FhlA8MHKBwAfDslxLxCiQcOaR++
UVc7qFRvSAw12kpGv9SiLvyEF1umsrnSf0Dacg9nE/6d9CsH82Zoeg3ecpxfaLdaTUAfWt5zyCzR
DeKamZQxkNldqw89/Jx0aHm3p7qnaB3SdZbqlQuTjeNwmdpWBnHyPwWKEc2FHBwzSyfDU/i0/vvA
YwOkenRy8MOCwXla0V0kBiohtASSItwvqQ733bSen1v2TAbK4qvc+Oirew3YIXPmkiW+lADTSJ71
uP0bRiZQBAMX+CO0Pf12CFQb59/PfuJt9uEAb6IriP9/4dOpsuCbsrHK1sIku0N29oKA8ppPoQsw
79gS8FWLHa197qK/gJ/I/VfsTnLHNbbD53cj6sv6C+V9yRLbfhTmbk6BiBc7IRD4BW4a1WU4dpAk
BsgFQ8wwUesi07EenU16/7HnK/gDyWS3uTc9tYJHBEtjPx/1j6avlHswSxbgEnmUeROIihFQ5wNe
Ei2W46AJsyh14mF7D/uWXYcNR7F8KX4kBfA3wV+TwFz08Onpzj/+Nkpr3ecgj8F+fl/rtLFpfkIt
ndzxnTmxd1FVkikYlD21bMqGzflH8rVGH4mCHFhmrT+MEkhy48R5x/V1pvB6ze93HBzrQDKrqDMD
L93Aa1TkFY6Jntv1APo4o4G2zGTy37KvwA8gktaJ92pHS8lxmqEWS70tAdsxwhvZcu62u2GcuGLW
LmzqeW+Q3IY9OkXnDP9J+hmXaoAMNSZ9hyyY6EQZqZfVzFoJepcJyNZsUCkzLv1giH2JKSnMY8zN
ndKh4t1XzGV158flelQLZ7S8PP2N/Yc2vWcVddIA3Jomy5g99eD3boizfor3rwEjJiePJqriTzz2
Kpk/RwPC+paNsRIY51Pj/mazT9LSWH2yIo3t+y1fMaI1lNRBzmEOztH7hd/F20rPls/bjpSw+H0v
eUf4RTAFTyPOpMsk/etM+gazsaX6Ej2CdIKjOQJBk0sUq7LeiQ/YGrrfMrOloB971LXI+wuYscAg
xH1koioF6sHHfiTAcTnQQui7+jHQNbykwKmC2Tyt4d5C7p91kEvZxghVprPFqxfFNorVTDEgO2MR
0LBsp1bOKZBeWTiJiuCplRlEVyGDNh5a1wJ2cGMLQbLWFNNp+gvvoHuaCEyYfanL63zoqb4TFCdO
emaoaCcimp7NVtm6ndVc6crmQ45SGZAsea4T17MElS6Wxh1Pn4Fmm6WdiRs8S4Txd2H+QmXyac52
hNOqr/4XHMpZoc5do3ltBTp/Gu3gr7hg+yLwqfAplqZ2+3UjFJ4iup6Jnu2X3OMYddf3+j5+vpem
VrNeRAPWEMXDAG7INXV+s7QL2M3EGseqJfzFkYDCHcqmkDK7RnvmmIP+X60gWKIpMzKCKCG6myEJ
DMVtbo2aBu9iKdug8j1Gt0KMbQWUpaJQYs2MBSRBJU+aZ6nVuUE53iEm270ZD0lEZWCNKbhlBZvJ
t6hJOwNpKFWtYP4khS3Df7B+777TkyK1eZ1Ju7EZsZpEDzmeWy0+uRmpM3xspvelRE1fNfwJt89i
IwiAeOrp47KNHsr5izDWXiNZReTV5rW4M++x2fxUHShLsUYsqp53bKWazE/bUcDotyK6IQS2ke95
hreBE2Y8AUQsnhFdYPxzH4QqWUetZhgQxB+hgVYQC7Z2DmiTv4SxLGL4xhSZC5I61LeQMVbdNO65
LkBt2Y+P4W9s7CM199cvKEwKKdL+I/Q/Dh1fcvbBc785gNhqvHkrIj4iZSOh0V8KiMdnmXG9lrr9
quCT2Skod/MxGbjqHsWyL68I5iBbIbHDBVXkCkWw0uHUt0kXAZbjgVALCWyLEXh8leccDeNvLRg+
gh8LUl2Ud7TPq1/cRuCMMNJX+O1riqpUNb2cF6r9EtnlduFyHecgbnMD4tQqgQ8/37MrKnVg2Bb5
bgJ02X6w4SXcLt3rPK8Au3Fr36bgcdE5zJi/GDKRIbi94zbfzNzC0purAGDriFVWaSKT/noQPvQu
EjTFNyZBST0/MybWEHHk349zu/SlABzN0d2C91GaUrEf+N9WEXGsLT3f/JlZk0DR7murC8g5ARou
XnzYos50ldKjUZAGU9Y7SD0Q8astxmssQ3HJDzcU8RW0/+8KQ3cAJ4E5dqUTZBsna3VUUSyjqVik
gdFS7geC5jwrNiXiyus5IrqE1gVNm0aK7OcAcCD5Mmz/uto0Sj/DTVffgyYzl943xZM345Uw1J0f
3elJeOb7yp7dxQ4Eng7oM4kWPZUupSdBfUdXZR/OnAnNoIzOM1GgEJFlo2IO3XBPaXm5nqHg0Pd+
RfTuNrLGqP6zOaucv0YP6OIS15bbYSLfb7YBRQS/cX8+UTzHNJpoPiVy/cbqeSSyQzsmAVNvOmcH
4FwMjO9vZJH+BYAPF1g26ewvY0zLWBLnoXUJBopmho0HAQ+ogbTCoKdig4grEwGH8CuFYMbT61XY
m7+SIQ7ta+VzZx/cP8Ki2muTngSZtgl72mxjjMxvXWiD6ZY8+kzplUN7U7ZW2yzQkwmFSDY7n/L4
ljUZ8ZCDtlIX11CjO6wtpJU5RO60DzXraAFqxEyzVNnHQm/0/000gkdiIgx5lwompTzasQXtjF+i
MnNpfXBmHGqvYxJSHgAp4W9LedcFxWw3F4A3Fqtevb7+wTeROHDIAE6VCC5QyyGZHdvvFCt7+1NP
rUo8hEDLqdVCFwlGAKsNvico5gUW31WHbu4jZoUrWtmkab0VWN76ChxBj+729nH9/ONRy1Agpsvs
LZdzjctF0CQ5iMaS7n/d2l1vbEtaZPUcqOq0fFYjD7UcamxoWyc16WfmqWNnvCh2UG3iFudp8rqJ
4mbBPzdHD81aIT2+IUDc93+b2E3GeuBB2+qSyGUiQLP1zhscEB0KRaDwyV4TtDyBm3GlQeCDbhld
XIcnnH0+usc83r3d2HSRV4qRSsjqUsV4hTdyQc2O+dys6Qxk4SaxS0bbj0k3/29CuSHFb+H8Gx61
tuHmz5/hIDjmV/49RKYJ8rqejWpFjL+WS8193toWFPdlGgyZlRhAUNc5hclVGGIawI5nrMFpHtjN
pDrwSbT9ZfNIThbFE4mreDCVbyJ1HjoCY0R8dDm5huWc8lu1tAEMVDZVBBCMupsIHdRlksqQoI+i
GxHmg2hySsnI/LGkgTL7YPd1PrPcT7l6e7lep4Fhad0En+tKWIcM0uk56Lso+BmiJ1XFFwL5SBES
0D9dY9dIfEKOt+qjxQmEek+aNBLXabXjXU2ZTQEDkLpuzRN+wEvkLNznV7c46hAJQHNiZhJvvWfM
N8YYYIjz9FIrYddgIBOgQw4Ov5UchEH8C64XmHywWOxdF+4zqmEapNeIpeX/TDiYNIG9MFt6gP8Y
nzEWB4bSzWNYoyinVdFotHc0ab5Ll6LqSlUZpT5jVde8M0viucg+33p6DykQQIg7gZn6lheOT8K8
hjjPUvQh1Xc+Lcm8pPVsfdUyoup2M0Ko7MGo3/Hvoh513l6u74h4rsmN6mQA//ogVIDyd+NUWefd
NSYDQEnrYuEHzBPhiU1boTWsCnm9TuDztt5xtbeGKQ6Of5oa83s2emAq98ziU0/axYiJoZgYFE8K
Owgf52ZSqy1y2TQoLcu/1NYhK+DTdslBPbkhWBh3Xr11QgVjA8uUN1uQuRlsRYmRRoJppAYLxKU2
nU/GJSmHCA3mNr+j1/fNUvtDsyXxkgIF4lBDq/c2pgsajIpHJKBKnirh/2B3ct7s7H8FIPzpkqgE
P4ZXicXvvaIXEiotJnHNQPfaYkuiUxEJTF08nI2HwAH6QCOGQt6MnkDCYi4G4b19ognRwJyMuaDK
KmPk8lZvU8Rb/Dgzd8jZQoorJ7hB9MOAf405nyPg2HGFVTEDDbdy38ttn6zTzXjk473bPiHyoNDV
wClhC97gYHpaa82zVpoa1z8PZ3nH1VHOLJhr2BrgRR2OQBzeSWwsFB7I4bXxO7vwmFXLC41UpjUa
7LCT7N8ZSKpQdBoPPyRPk2W86s4TK+7zmKOKWQZXHRJ6rxSroT4k6ROdEX2RGBfKYBzvVx6qZ3aS
X+R8CPEvQN45p2KJrB0vG/9CLYkzmf8ZtU+bkUPrJYvLFXMYDhA3gLWbLc7w6q0yxlXNPKtSp7hn
+wp2YGoChH9wcjpTNDeKOH1EjOOmD0Gyh9MAN8QatlDD0MUR9ATHlPtnkBaAQwMQuhnF2JXsdTxH
DTJH7F5QZjhd8iatublUyJJ8lG37QyPgGF1aDXNP4eVH7fFl/nF5ZAznWvVAVI1Ys/fsz8EWotTr
pcxAS1koOEo6SFqchptzeppnK5GuFrZoKxHVY5wVLBAFgJOqETx6/SXfkDjSB8Xgy6ERqSaYiRAx
et2hjnGuvtLKRy2yJPCwzTBhBKIjkOndI7dqDAqzVF1odagapy/m0w91PYeDwKboo/U19MShtf9t
Z10+rO1Lw4gue3r329WdjM5wUaF8YRFQABrQ0WOzlZKYMQjKlhOvYj5dAJljNMk27P29ZHhbR+Ge
gDdJ197a0ux76Crx93GlVmpZs4Kfdv7kmWqxCk6Vv8pm8Q3mY0neV5mDAusdL1wozvYZxCo1/keK
02tXDksUaZrHIs15UQU/efjD/RxG5+Wk5qd2BBpodHb1zRko2AHcVNv+7GG1qSsblnaTRl4EN7Ms
Wky222A2/Jh2L4N7BaDvbP5DLGVaOw832c7aMYbRExMCJxLrZ2LP6+ppv7oJFh52Gn+iN5gcmRqq
cQpNuTurnTjMA6+4TgdeMrb9t27cv6PBRVmqUoiw++FAuea13p2s/+tORreUNdWD0jHGp4+m/qRh
BfCKignsr/Wf2dLD8zAFi/O4YJqL2B/BxJ9+b1LmFrWsqcAqHWtLELidq2REsYTf74OQu5m1CA96
1A0Kf/kh2CuI4RntH4wwlZPqIN/X2wwerT6Fv6lLDh2J85J6e2b/tCoC+K8jb17eEmHEtFUbc3lG
/igKFbq+WzmrQDmPkuaXsKH5jn5RmGMqNPtpIPmWh3paDcwefdhwVZ5M+bVt17hOBE4jx4eqMZtc
URm5L/4i31Q/TsLuVQdR+WK5DP8a4Z7fy9ZdKsE57ctwSheMcvRSrzMA0ei/pdDC9Ctm5ARRmtOU
2fySxm6uU67ykP4K1u3lbxgxpYjgQ8nPRVPjibmUpT+iqAm3Rd0CydMhImylYFB3rA47RVmJwuMc
lKGv3ViHCmwhR1Xw9BS17QYSvxx9m4VsCUJICFKZDL7nHfbt/FHcZ88NsYzra5OJMuNm8Fzn1KZN
t5vEsCE4nCkxqB8AkXHvGzd8C8eSGQnBM9Ku1rWrQY6+VuHZMJex1SpsLuZ87oQYgb2nYASTqE5Z
nLdhEi3ToVfSFGaKkCRGBSjnAgHETZ3+8QgI6MhyLoUn6G4LM01N/y0Jq2ViGYl6CAdwwXRVsBz/
ZUuSfeUUlu+ECeTom4M/hAKvZo08gctL9hT30ETudaXwpU9OWqdPtr+0F+61h5TjKl9B40JjWyHs
G49Z0ZOAmfuwD+xvRRdgpmDijJmAVe0/xPeaSK8RJCcCJXExFekpNMNUmBS9nlzrcxkNLxeeTQba
1UGTEZuui70aV5GGXmKPJ6CuXhKEimhYaePJoAZuYvAhKZJb8/goLOCDz+QB8NRTbMvXiINmFVzs
0X12To45i/uuGXGPcJJmfhDt9KtoYehvBXnaTQcOCOhnKfCKLjcSpLg5CtkcU6ip9Wd/xfZavCvZ
XrnCGtceNBuSEs4UCURPbBcwp0iNh6Z/x4zrDECrGqO9WY7LciKOY12NADxOHTUXNOPrC4rseNSF
132euW8dZIYRjSAKJBWbxgR48XunQTKSNzCPyYnC9FzGAND0LJ+a5nsv1C9PuOBcix7sj4yqO/7Z
F20m5vKcJCSSIaDWGUTZ0Qcv2Y1Nn7E+/3ROPGQea3pAkstgcd1fCqLdAdMtMT16BLfSYVnIofk8
pZMOJaPPf86oVEGjUCkWKKMyTW4H+gcGghAOlycFXP1+EdVjwjgui/0eBY1N/fEK/dxXGqZdPniu
diKLDV77WwSEecb38S3YAy4a/j1jtI1blqEnILs83HHXiS8VjuZ6a4xuYXk4slpScqq5SnQwHjdA
JQaFdPZ+W0UMmrjowUG/5FqvPl08ZviXBbmDdZx6YPuT0M71o1pxr8WKyndWiud/28m+/BJWlWj5
u2bYpq8gH47evXbpnDhwQRZ/3SkNUbjNV+LRc0S3tWWcGJO8yS5kbU+UiPJzFWpM5nzPPJ7a0dxw
w4pzQlNMmt4uKEOJ9J0PL3MT2GlsjcFK5EVW5+8CEIYMe3lOT2Jtc9PaEdjPiDqjt7Y6aP0AUy0n
wocE3g4jxCQVJw+qpbRz12YeBB5zpAlrzQC2//4l4KhDEAn+vjDxXbeFCYVm9zGRRb5z7DcGgOha
9Zh5dR7BzabVIEM/HuncM6P6hwjTqC+lv7HI4LBUaq+Bags05EEoJzuvBDf/9D8jstJQH0pw0kyr
mGwBuR6J0h9oOlDz+Kulm286bwv83nPdL7yKhWDoDp6frgXze/r4xF+jOmmlQyB2eB/IdT/oaKJK
8KG/4KTzge7r5EtuKMPagcVRzfG1MXQtMHNX03jhT6ESVfyOWtlAxzDtZkYSA3B3JuxGT+8tIX2S
MjE8kUu75Tn54RIl7bpTcJPq3He/zF4gyrLGoA8Ev+IfUGnI2B/QsxCX4qpMCA2BRXrF/QwgrgOf
GbAs3ojyT+dsevsB2V6NYUkDfIJNWEqwBx8Gu3LqoPNjswsncabbjCpHEnWA6O2Eo/g/0xfazia/
zf0c6PKs78OlUCk9zsI54diPYOfpuqe0cnto5l22AMNCWNk3dYyhEmM+1jGurQZIXZb0eVL/N5I/
ENgbxG9o4p/VHuS6uMLzY3sJ+fLnwd9Cz0tTF6B4mLl8ITBwDCQiyTlypgs7rm7XWSogeIXwLTGC
SEkzjFCXpomfitjzxHBUWDhWDVUgiHHNm7uV637SUztG2g+H6+PSCcXKRn66SBzqZc52yRaTvPJ/
Y1xCaDW8zd++9HBTI1p9yrnIdOteLF0lRpagCiMi30tD6pDouqlhnog/4efHM+V+jBBWV1m9YJR9
0I5svIoSrNbCiSrCw5iwhGlG+Fpf/yGvvV4NIWMQu004gfm/CnadLfEJcIrzxoq8jpytN5B75O0C
s65I8JC4D5GZbmvKyitZ0CwtVUsNEqLw5SHQ/iqKRVLJb/Ok2inEm/ck02ioO3HjipuZFNT/0YBV
nU7UzEC3ltvHgSSmWh5NMBUg1bc1XZ5/xrCdZsbUPvFR63l/2mu3GHsHFHKkq0ahBraDQ/OI66N/
5TdLyvjK2M9zuX35DsGly2mM8WG8jXfP4dyAyi1B5nFeJqRRcHXxTLPOEU/OsFoolbAfHLUfokXN
JZssyUVzyD1//WBZbcusqw0IsNqT8tF+KS7hLpv69+hCqDrDtJScPVfDhMamtXXjtfFa0I3zeQUt
LvtKBTGnW5WVMBmlw42OE3+weHFRyB+yFkqNaGOqvRMToHkUu5jjpO4RDudy4HqYOcxI7smFJawN
q5mr1dBlV27R11ZdPD5HRjLW1UZU4hPlX9Ewe/vWzQHzRcu09pGtP9q91A12yB4OiWHpzKO0thuf
rcSk3y8ygDo9U4pztj70Hf3s0N3oswwP8O2xpNcetTzGaYZIXDJQ6hTs3QtITb66o4NwC/XGiMfC
xbs35bUNgXwmICZgejyNVEf9iZugq499QxBRjEaaa4yR8qC0MeyQanDqF11TTiVCqZbqSnauTe0k
cxypRFAMQkMk6jH+Eh+HULg3oUGAjbN0lgmxMdU43h4zjREs1rfQBG606lw3TvSeFpATFrJagDju
SU2XrdWjZHZFZzkrmguCF78T1gYiKpxnOoPoAUDv83aot6Mw1bNEWv3JEaOIaBdDuLLXXYFc0pJ8
4Oo+uzDN69PATEau3bXJtT7cD8x6WbBeJO2KxtrTgPri47L1BZDaIHzNkRDO2WY2HApRmS4EV80U
VkxjIGM3myC8ByhPm9di8dK2mMOZrLfzEPa7WdWwCjIzZA2j95lrcvtzqRbXSla8oruqWnm2DqJr
MBEhkY+AedyiRazNJ+XkL8GCI/9xOixB52ZG2L3xR0XJNkPIZdacc9EBx+dgI9uBXWEn188wvCpm
wC71x0YPMw0yFv59CCFhEr5Y4A0t7kzfgrgDmMXx/wO2agYEAGsO6mQhRgphUCtUxhEMasfDr8nC
+/xjOuOFNfK1fao7+BbS7fQtjpI8kh2yBt21Q8OiDM+mNSFgiQNFLZGV1TAaL5okWLYZRcIoavi6
EqSG3vSyJl62glz1U+J3Aeg1HcHQgjmkyBlxCrp2k7hzoNZaMi4Cf+/sKKOoedtomdpfxlpk2TgD
cxA5gLnltK+QiVYCftK5lzGMvgGeVFZ/BNYjmq0PgTjUvp+l/3qXwenrxGeDNH36SK5buUzxrvKI
o+iF5OR/lso9b1046BMXPCmva2b9bjmkZGG9wrRy69cogFUkN2J4dBx+rw15rnzzXT8sVYmpkXbN
+gE9rh94Rril9M+vsMpE7Ow+zG750TCUNs+C7jjNjl7StcgZLCgQqLxU5smAyqh1z9dlmZCrYn+X
+Fe9yF9DnOHTnxDf9VVMCcrlPYHhQKhYNkKmYwe2uE+OTBciJdsqaM/ivO76gEetgnAKtFtsDkpZ
/slQBLzwBKETHssrqYaApDAKvA27pbNho6yijjCgJSSm5GuqFTcqKTe5VQWfxpdEdEtkYmhk2r/a
HOz0PCytRm2pwuoyKf+CkANg5UDVDx/NLIm2WAyeI0TnXMtvVCo3nPjfjqjAkCT5hb0hQqixjIAp
bi5L8hDhxuJxdjTck6hGhbPY97BgtA6ihWVs0oU/WwIvaq1/b2h3GiMu9pOcqMBfdBsure5Gjw2z
hiM9Pf/LDk1Met6nV+uk3ro8+po++bHrfRpLW1NSMjDIXuyGAxkXylfU/0Z9ruGCiEbZLho+1HXn
WwPH0RIgNeNTBMY7jRgrMqPCtw6UoTe5HZPmAx46m4GdnTheuWuYYhKz6/leZV+CY2ua/DelUFxU
Z25Mpf6RTLb9G+4AQDMmUmu+zLGgRgkP9P5R3DUFRzQkr7yYR26IW/euPtlKZkDL7GfqczgQ+dS2
FAOAjU5NttXD1zqDyJ7a1SFUpfutdUz1IInE5DUdDgQjtTgZXdSs2A6NMuvMJgfNyXEa+rdgno0d
BJWilwgTJLjzhqF/OgiOV/rKXScyG4p4VLuTTK4ETQPzcFgiFQTrVrylwoFknBZGO4DyBXFHdihx
ZIJKkOu1AoQpa1XIe53fDoGYxsbDVgpw5/vYg/3UEjE/QgywtQe4n7Jo7SLemEg12wJvoHq+pTDi
MN5tDKB4kyVAQs9opW9m+MdtVn/v8HkzbaIvkV5g0GmbDogp/9W6H/BHI5NG2Ubb2+h1Zf/EKoZh
ry/y+ItCDQMZolpFHYJPWCChOWj3WlOLtSqbvuqOG/Wbd+vmlcWI7I2uWeXDJz8QRf2MWo9wqvcK
MvRoZT2mrmttWBZYTOIgi51oojGwlFvxROlzZ+tk8COGNy+clgx9G+k+gnZoXG/wwrC9Lcs12Vib
KQPdP80YIPUGScKl0E7vFpcCVepaM6p1lEbRQMkfrgLeeLonz7HOvEUH+yPDBaAPvAb0EmuX5KKW
QKZGnZsDaW6wNiK0QtIUoAnBG5iv2BgsZ9KS/aHrZUCpPfmLFU6At2u0cvF1awxJo6j5rbKbE/nt
hSsmBmRfkTwjI1PNwdnVxTfGn41eCw1BjfwUOrYvIAs8GPY0LBv/Tu4FbxrDRlapwslU3RX5KgSV
d0roQxfUO9k340O0zEScU3eAKsIkTj7BfKh1k6kHn8Jw8D8aOMjK0pU+8fK4neuWkKuOj8mEW6Ri
fsbfIedGA0AQOZfHchpO3tTY/ZeGRI9VKFsMeA8u+ioYmVyDdmOJwik1pVN9FC3uDJf2kyc/bhP6
1bts7CComr6xIVdMGuUkw80YShVf6j8iurn0j1D2irhYxBYQL2UH3jGfPJbncvmNumlnULmZpEUS
TAdY6N95oZK1tVJz2gOWHTkyJtMgHOoB/udlKXFKyJYyzGfcA8vGwlR359gje1xtQbMEkswHzzZ4
Jottb6iysz/9csWIEvK1plU83qVbo6+apMwPULXBUvl7bSdK25sRqmDLiQOO1yF0YwJC7crxcWQ/
2TMSApMjNUSu47Voe9Of2tQdTJ/P3oUkAUbH6eeToSXNXHvk1SzACilYvOvJYLbIE776d37ea4J+
98azBszmKMdSQZoEBDjNziyvWfnRaCFdjPhFR31FJt4lslYJc/UZ0//9ROLLfEmMVdPyl7Py4LlK
ob3Z1DOoaGovvaKROvagNLZEWgt7Dfyim5TBsTdt3MOOz4i1psBoo5WBEZfrxklCuSayoRShRq/6
QerCphWj5OnqGBON9ySadoAfsI/xC9B0XLqphKlABbuHdR2jIZu12IGVc7hIztc/GWMG+UVXtbU5
nYMPoBPGd+81uoLcMzTiptwLH+HgQcCNZ4u/hD/TOvqbaSN75lFqZeAb5GAG6kFF+OVxEBOrfQ09
fjCpD0qbgJgBCXLatQlYXP5533DEcZG2T8lxwNMXCMh4DtVzAiO/i7CQNjXL6p14zEYqt9v5gOpF
YRuP+g400ywT/32CTqz3pL8g0+WP+8uZkp9P0g9ziJQbU/wEwRKpTWMW0cmoNR0uACmjTmxUNgyt
re+prmF+z9QADKktfwKAqiBPSZQoqwRka4Dz1KOAZxerc9qVICBQp0Fc9F7fjuOf9CzA7Epia4n/
MnMOoCoBs9xMfVEp23oT3Zq9qkIOT3QMn/tq6unlyYMp2LuUZwteAMIPhDOqTNYx61fIoImOwXdQ
XaXqb4gYTbMR0y0QWOHhH4W9qush3asB2To9BsdBYeRIkR17yoj3YxcJB8byT7HqgoP9cFA3gbZl
yEetNHPQqL6l0BcLYEt74LQ8Na6wUx77Z0mTDIjS2PhZUPeRK0U58cRcbRoSjBD7P22RaNA9IYcK
uvYKaQjYPnVJHdwg8LrKmr7yyRQUgJdH/g4U4LUYsddurcEDls6CRRIoSQIUnzJxHerMWAc2g161
5hLCD8JiQbEVdXqNNCNYPEWa6sdmatwLKJAn24iKzW/Ds0DPOnGGcSpES+ep93txGWZTdU9Aw734
IvfvDGymuMkCtqBO8J/CF369V3kRIawEwvqaZ0gpn8kA24fY7ygoVI37pXNdSwAoShV3E1fhBO08
IXd10ydZEb7N89zFQa/GyKNs60cLwI0xJd/GOCkWgimTIdBAtS4v4t/9Zs97bzM6PaMier7mujeP
58RWf1fHEDTxrPxhTsEDrafH5G5UxhiQ5RhwJGGdSnnt3sJbXwNR8fxDU1PPkNIjCiwY+TYghIL+
u5gkOqeU8yE2e3sH8aOCFlnyJoRQnkNKMxOFCXB/BLN2lx/A3b1E7iS2yo5Nqvi6+NcodynFqVwF
E8nUcPUOTc/EcV1Xcn8oXN2fV3tC7VodQahw3NbFuF7TSYm48RXKbzCcmldo6lDAoerKGsI1cSNs
iJEsIOOojZnIg45GZLA38hET/hTPzoXzUCBfl2o9QkTyY7owHyEhCMoaQPnUgdPorGEDm7kgY6VJ
TQhAVyuk5aEdnWkLAA13BizwYv3dDv+5y86VqSj2TGsBjhsMsl4bTi5WPjbsxq1EMVamTHdxPpeA
b/atB5gZSGp/ZEQMRsZTEh0V8W0LxSYa0CWtArZPMAX4tZ4U3W7PLh43E07rtthJ85icNfU6C6b1
AQpvsIR7E46nojCXIaNQ0hK1FmGg9qKWkq6ZBY/xOwmEaC7S8NvXev5RUPedfib0j1gbfRuSaXBT
wd8Ly0kidiyZRaImnszZDjF85z+rFxDryko86mdoRBE2S6pg8eU2z2I6iQr1CEGOp9BQYq/WWj2l
T4vbBzlZCPRqHC6wllERY8mCWgPIzgX9CvF9wAxAGYP8N/TfffWXAjqeXWnmIKku2iNCWTvHvkpI
mW41r5y1AcQk2huATs8wPtVDF23r0X8wViDl5nk1qohRxzpZy4hhu7O0xWOynHa96lMbAohHfnKI
Fea73+WxavH96IisyjYNu6fETFIQLW9ZylZbv6N2oobt0d09+edAqG4uqVNkSNvRTCV5ndd+BcWj
Ls0IwEeNmvwysw5G9YKOnbCXh6OMs6eudsWLT1zlm3m431b+ZHimb/Q9ef1nZVvoJyFxBoquZEUz
tCYK5QKeqRZXMblOj5vWfu35CnyoH3QT+iuKQMF1+mGMMaQmHOSQfgn1RYVMEwYi0ZmCi0QIk8EL
W6Uilc2m8f03SpSVc/K3zhEttOsDxIeIheQlBSGTNPiwuiS3P7bYtyPfUTlnmqPoWFGf7qcNnewe
0EgFVyUsogLQxWj/Smsjll3QirY6HWfcunej7yNLXpounOY2zRVW6SeGI6bMJObBW4tMFBHbAhoA
HeSPSZ/Rw/b1cIt+/gNy9cbcdhczmPVJuL6ClHR9j/7mEDNlCVLfmpPGX6appDQNxZGwdaLij0xi
JCbuSy4y4pw4Pk0mAiHer2ontlF++1EOmkyKq4Fp/kBi3vMUUKzTRun7/aiEOc5ZKvWhYYsVk/jG
153hIk8qOtVSx68EN+rBnJk0uIhQkiI4c534600h5bM4IA5oOsr5Ipu5tgeOxuz4vEokzChHArxB
cosjCb5OYpgpqkZt8EBaln52VGiDrvyz9bwyJMwWX982l++VUrzmwImw961I+VQpP/ri12ku8Qi3
BUL30RP62lbUDoFTOgSyBk+Cytrqp24MHED8O706IdJ1t6GgB6KGCeg+hn5lUsjZYM/5HLk/Aa0P
wqBRkdYg1PGEinzIoq4bclOcIhkTQkQEtG6PlOa1Z2PHk+tOjbQLJJVjcosndK+57CoerdzVcyDJ
GL3ZKmbKs4eIofrZJyqBPNx+CdDlCkNIdZI9qSqjOs8e9isOqZBBuktVfsKtH6X3rAj0V6hMkS4F
c6PRi9035RF5WYhY7vRaGh+d82SFJJQIcRX+cKxxJETmjoQ/H8ekGWZCgwEw8ZqGJbwfSUCW4v3j
K9Lymhu2MIOK0EoBMYDN8JE7XzP5MAC1PHBwqwTO08qk/pl6FYxOYU1wQo/ta52ITTnTkRhMgzmB
JOYLhoEOd6D7ZrFlFeINwZTDuCMmeuWbEa5V0ZmmnyaATrk/Q5X92I0siE4dbIVE1D9Tj5bUv+VF
3FAROR2K+15Ybwv6ZSh/CmM+6FC0mfn6aLwNUHLGOdlijXBuD2mZ+TGVgDXhULek9UlBH93RN2FQ
f+D679abbpuc+g9Guj0QcQFD61SvwFAxSeI6p9jQCogAPUgUfrj7DIrlMfwZ9ZQKi3GT6piPrG1c
76C4Ks8LLxs64nUpJbSjIyX/eWUkx5wpQkWAMph5zDSj+MEKkMOdbPUi1hnDNXafW8vHd4Udclox
jTo0WajoR6SWFK29Kv45Cx8So5051lLL0feObLX/A7kb9vcr/VCIHcfaFKrnLVePEUyjp3O7k4ES
984J6o2LwomjKAa5wmuIuQ9ycPZLaijXJmwtM4LXJ/00HuTB3VtADUF/3QP5Nza9xng7vjeIMLbd
08pnbzjYOnl0AlkMGNZKBvnUVqGqRXOYNJp0brvKjDvH51qPLH04J4lH8bckkNJts6zLH6NxFx07
yNU0552EJRDL/3hLNT61L7HB82jwBAECIpym2xpu7r8W7ZN13TdrbgDl4KUOpn45sctqWydVgjog
krzTEUB5AvaiXJtgJto/oUNlpoIIgwcF3T/DEg54F37sWuvQDZ0wtHOwhJGqxHBUluK0ETGFO/Yp
6heiG06/xAKUoPjvFJLCIHi/eswjef89E9JuwJUMIssoQL/ZztX8tCFDww4jZ5ihZh9G1Hl+1nP9
zfs0m08N2xvPi5yJXOV4BtSn6BrLf9aaKGPDg7iiUBIwev1CMe0WYLkEgAqacy9KFv+jmmR4AM2P
jzhdGNvRGuKSV3eAfcelIZAtjk443pTFLvtsA/HIazDiNA3TZZr66+RD9zipNTypCyxp4alrQUDB
HV0cBYqm4LqPPUZvBF2lYjDuTfYSoJKM2NBQnNapJ93lxLaKHMJY8pp6wHMQo+kHBGrNz9X/usl7
dWFQpv8/XXe4O5JKZDDYmtSZ/uz0umS/L3P6AQpMaXI46OKEIWrYlfXxasTFDy52TS9Zdqrduavj
TKokel7mXVeJ9KX0Gtj8S8ZfMT/7TksZZ4PZ4OMdjA9nHGVjj+LSWDacHEW/8KGpmaYGHubehuxc
nAzmHGFSl3DS8cDrrAyqU5MLsOojoVp7J6X8yg3RWc92ee1bwns/iznFZHGxYNvTNq+5XWMr9ywA
Nw1dd0eQnyhkWc8+I+Rr6iEdHcjIEMpTH4W9B/77DEmwN80QwPkifXx6dV3BMAgUCdmwYkkIe1gX
r390MqA5M2vkepaA7dZLeUfWD31d0sLWVKB2XyhT71utypEww4bTaR/uFufnO1sTHVQRcE1DWFmy
ot3UaOHErIMlOIbTnsZ5lGHVB5j5MiQ9VgkdSsykwfPYnW6CtQhS7t7lqlkTXlfmwlJL3gtlDFuU
DzZQ08lY2abPtp0EnUnK0OGkStiFHulmfdUTYK2yS+vs2h4S/wL8eQ5NPLMgd2J09cVHZH4JfXim
NmaTMuOifqP1bbjXqyMJ5TyL/4QZCbWiwz5cJqieB0jKl1ziKGmDcTsw3lORhQYrprjNBGaQf325
AvgApDNnQPg79I/5D7Mimj1qS8k4E8UxJPGJ9nyiSKBxIXgoFCEcJkFvVNjfK5X21kP9sVgH0UVF
jgZA5TuI5immfAfT50TJ/OceKGgESyOdd6K0ZW7vODcI48X9eW+vBq9sb+ePFh9Ykm2QsMQIv7ci
XwiILbos0pDkZIUbPzTEXtcyvMTgAmL3/UxXmdCuCurwNpmqpMyEUEWEV5hjYoDCTwvdF7Lawbdu
G99lTHn1xf/nw4kNkhbCnNE0GNiRFFcD2VpSNuzCnOgxiFLQvGf+BrCMl3ByTA+g5qGf1swHvEri
sOkTs2CCVCxnVe+wD18K8ZBLIMK9QYTPjmpETd7Pwfui167weEuKNXZRKD+CIS9dB+TQJU1aJeLU
AA41Ou0X+3YH41OrjXq6wDUyHj9vIrbA+huRX+HZiHrcp+I2cgGddKU/Zmwd1VmhNZYi+9x9GyZL
sweHJ4TlJ+meJFFbNvWMVC7IA8bkr10dUkdrT+xQknsbnrH4uKQrTv5yIRb0s9Fc50Q7S3dX7gsp
0ZheLRikrjIDgA9gW7HbC0fV1s7sboszcX1IfBAjBREOLncZOh71WFaKQEtzpj+FUbSn716I7aPd
zWn4ls7vbCUVJVQu3/5emwFLIWxPn2O6LW2Lt/SRqpwkCgmAeo9ZbEsHGva9G+pAxLLfzWtaRHIn
ps1t01UX2oUdLaAreaIsY6HWlYWEDhuRElWogyZ2eJUGMsYA90SGF0zH39xfokYmA3F55heVtRsj
lGPnWpSTRdBrj5EEYaz+wqlg14PGWfUEvJy7cjkv0hJuiywQTwd7U76e8fGtGS4eubkotvgtkiYP
frjMyVPPYEour+wbLGnS2vkA43NJFM2Q5UEVbuupUxEfmaBWuVx9iQiRPkpK22OZIBzUJ+weLtO2
nD91IEsgfOEuAhveWFzyE51Rx4VDLI3KTOFo7AR0djlYSP+e7YJkYQGA3lLtw+l+ea8C5DQ+saC4
vqbuRMfu68KTu/J0NlookRcgsp4ay9ludTrzeMxAIdFaQ9MWdE7fovI0lKi63HjYmYMOGODLbfpL
igPDLfWPF4Klv13SRaFYBpsRgva2COJxya0DdJiX2Y+77eAtXyGLHDAJLnYebbfnZS93hxgWCUHM
w/EcE7kQ41Am8M5iCQHAjQhIhU84dUAVq5x3k2C9FTzkeF2ttXWVNrfJd4IvRqfCwQBwlJhOGNJ7
FDHE74JeH4kvfmkQsc0D1e57wUR96DPBQLZj5rIr8ymcydpsDVJpS541qBYzFC1YxDS5s+RO8QiQ
YPgTUJ7E02Qv7i+JW+rbwZzZ2MRhXXZ0gLaWzTTV4tMnAr7AvmpDAhQE83H2y7kHQ4LBlYeYeGsg
P/ExaLspo7Z9aIQ02bRfqn1/UQw4S57nDxxgdtweQKt0aPA8ppokeamh1jd+FzDJUKUEBP4a5V7C
aJPOP+PvZEUIhRTY8AKdd98XRgFY5J9eCFWVBzmCMMi8aE0FEC6r1f+trpywdwFG8PNkZw6sNLnd
FNrv/bS97YLJDbDww3yroPvlwLJcroxJGCqlpIsRnW7mwY4k7u3PDw+XyXBCFQ8r9+fIk8oStjq4
KjjYO116zf+NwW93Uni4WDVsK759kF5NNxEdZm4ii+MiWsgaeSGp2YnCH3oHhyBYii51rCo7YvNL
IbBLyMZpWvFlI6xpZAmBvrf3jImhnr301mOoiLNDSoQrnk8H1QDx8IbX1ZZWuKciM5iRQHbDM6u3
3ej8/OgYjUYnFlXhUvro6DJHD/El5cIArgg0Mq/e9/JXqVlq1UK/pyKxCaAdrtm7BSyXEMYQJwCm
oXsl8YsQSJhYvFPiqUJIM8DUP+fUAEideZ3n02giyhbWQeTU6FusKWZyyC7zNjQQLitu7CFqm8Wx
HTWpZFXXslKxIlf55nI5nRR5Aqwtr/Ho4v3AtYXoN7uQWjy+4Ck45DxCtL/OpNIuP2yq0eSoyGo2
li7cj/I1QKyPfsnEJOLYFum8EoREYnGYvtUtR5iEzoLIVDM60h0Aq3QNXRhswcHJ5S8b2hyOOdDK
yVJ1+UkNMCOeh00RnCgoIPDhf0ZIdH9QNDsI/zGJsfTY/IHZ2vdX+U6GCAJLzyJHu4LkV0sRqucc
zK/5GEATCFqaQHeUQsjx3Kx1/etiz1oAkaizWsPXiC4d7VgZ1FhrnDapDmNChBxnxe/SOhU1zACn
CPZmHS+sqlZE5ZpIKO3ErONbxQNM2Vek6TN2MuiuKGkQ4kUHy4rigsZoirQYyVxSh35NRqZ5CEAZ
sfv9IUkolTl0Zjs5BzFTCwoL5QkKAofBaXyFXkW++jZv63vkHnWt0irlhPFzjRvCvwxNyhs1RR1A
jx4tqoOuoYbALhcjB9GEb+atpGx3h8+5e12ajzvNoFH7Qa04hLFk9qZF+ExZasTJhrNxnEgPgs6j
VG/DBUbr7FibYjjevhPQ2UGkF3ORduTRB6AFcWYdttWE2J9K9dPuOZQNlktj0N31zQ9NjsMScaQK
FC+sUOQI4fO32qkFRTUn+JMKfxnTAokIDj54IHJcK+WwfZa99bJHtUuKQ2ML+V7vTA+qTva5ifdY
PUg5Ws8xcv+PHc2MzZq2U3/H3m4u3hMsk4/zwOSdk6eEDXcQ5854x7VI5j+bFMXnTIX5kDp5h4H3
VA89ZGakEZUDeDEsZ9JYPHKN/BHLAgX96sjTcUkxJikFHmfiXykxIqdVzmAjCLWJTZl+U6uYXKwt
mCF21Y9TObt0Bw9Jt+CxCzX8CLtB0QWO4qYKnngjHvxj2p8qtz1ceD9CBlcrYbj5T5Cs5oyJ07/q
9AsUNYn68uq6U2ag/qKmqkh3Pj1KsSfnxhBt1NV/WRrAC6yq4ALhTMBZb4yuMV1VzrhFjV3RvItp
iKlPMjAvdWCpYKJ1CkPv7WIxYYBgrylUgXGc8YMDbBPRLDu5Qz+JlKaylONCjO5U77amfyFDWicv
CcRAEg/DznoZ2f8ZESe+mTVdHxO7xR/xfau8miaIRaKQbta9zr5ucDaYYubR2qzGpJ1VH+DaChRc
VFs2CCrY4cIi+utirwi7PJHrH1q6nFwNwqtgX21wivefRze0tBLE44h6lO4uwFKcJd2/LBrJEdxZ
Mjd7Gch4wOqxhWF3zRyTms28GGbf5ElINtv+0PRDHFfxAILMVCfep5ZPP3EBUx+5oft9myilggIZ
TcvqLRYwaWwbkgS5LOnKlAOd3CE0Rrw5YZR1Fv52VtWi3pVeCRtFAO4bjJqmC3p+D2CWKfeq867A
980bAN0JIzNXFtRu3al0bKjGk156hNRhygkOL4bOOdRFV7WmEwWqhK8gx1wR5XNvIixpBgCk2Xwn
rgeA9ooGNvxEH2EF+c+FbF2TsI7qltdxpQ9g0qp86DKHalm9jxNOXfC3E4+VjyX6NKcBSLogOD02
Ysfsad/5yWMpmW+y2lQqsJWTe0wlS88ziBeTBF49JgwLg9jGFJKtukKBa84KbjbJjfh5Z5ZXdxYX
pdM5E25r5YN4S7c7S2qLQCk0BLZheFhbO+m8z8ooLe4c+gbNLxWRChDtYyEglKAot5oI2gg6Nnix
0Ru/I1BDdVzgaEI0ZVsPuru4KhGlHNwC2981ISbeSKiw5kFHXpemiLvKuavQq6YSdFXwCVbM/Psl
THrQEnFZpXvSp3jnD5GY3K9MX2pkvLBpmlLabWksgp6xNvex8kPSgl03XRXKTJJRKFr4oRrZjeLT
Cy/mst3q5acZZzJcew2ctonK2rdNdgq0FB9GjDphr+naa3rKJtlB1CS1qFvdaN5YWivS6BEvILEr
4mGBcI9bdRFj5a4b8YMqBzNUsSHxGIWrGTbwp5WggPv7E/uj3iz59IbgTUtNx0mMT0IJmnF1u/NJ
hv7PU8dIn/FbojX8w0CqL6WvPzS1jKMZ0kWRnA7xKJ4Uo2oHl3so62yxJAFkTxxSuT5bFLb1bdCA
FMN0cbdXMNIg1KM90kV9RUT+K6gMLfkPJX+D154BMiuLjKErVgRsKjvUFJguGEyrivYGP9xS0u8s
qaKm4SX3LG+hiH8jbrepweTLJvYL63qtbC9nhO9y6zSdTOrdthisjjRMQxSWoLVlNfPka8upTD2P
zTWw0OH9Y5xKuQ/4Ju8V6irN5Q7jHHHy3qIx4xDD2j/FWr2rpF+BVyJtSdH/6fIqYkBqlX41xu87
W/rUCY/+4369XPN78y142z5Jg3kpvMbCLNMyCOe/gk9Bsqz6IkDGCWRlIN6JdC8WQUUWI5te7sIO
KCWKI54qo5Ozlt8xkPccVQ9TEEA3VJIbX30og8xJITRVn0OqiaDnKNX8coWUWnzQRfiNxD+6WQue
YS3kUI+6VIfBeo3nS2pom++rXZZ17IPah+AP/nlHNomhYTKjbPrzecHTy5pIDGuACJdAHB5jAcNl
/w/M6umLadpdIBE5e//vdohAuXHL8sbbDYG2XW1yfNC0Z8cEQbemG7BjBKHHAQcNeLw0U9h2/j3q
X63RGepWoWU3W4rPFsrq8mqIi6W5Ngz+OUcCecYj+/oGcLRtt3SFIa4dN5bAx91qC5uFCZy7Pi+H
ogC/9NxWfkWWL4Y+XpeodCtGzEl5n+30uK/Zc/twYlphqTpNbov5qNBiEQZpWHQgwY4lu6NenHOv
eUfo1BBtq3GpZtH3NEagaSQjYdVLaCNtynbKrWSbotC+5QTDawvjXNlm86Pq8lmicL4ErHYG/Zg8
XhqXCE+xbR+LgWxTWdMzWYv4hmiYbpa3OphDWUPRNejGq1nDd+Bh24KQlbUSLq2Vagsp4S8wAcH0
Ci2IMBGaf1NtAC0nOYvlx0thUpYZUl6PIyTqOzxHDC2Jp/aeeJ5PiBlA9PnSKcGUDMe7zyRsF4G/
eiqm/V5SsRq+Co3wTiHwprrLJQ+pKBPerPei3qRpK6+376WqFlOJh/WyItVrby4nccTo3Ghl8/Uz
sHhpqprX4T6CsPTNJBl7jAiYORVFU+rCEzW9kIoc5M5xYlWD3v/WZ09KKloI23y7YpUTuJZGXUci
gk8OO3gkfVtFnMif6dSk6b1DcQl9MZEAxTM0xINcR3j3X6YeMl8WLTm0tGT1FPvur5ZbqaHph9ZM
7vVSCMuWe3C2cA0dsVoxZlAlwNMcrooaF/BI6aPZnX0/i7QiY7fxZlOWXP371NxiwJDDLsvqsHWS
V7ybxqgP3egwtwetnIvLmn4ufHsdBUQHy7o8B0ySmumElvSNCqDqkAghf+jEXHAFlGiZMBuLoX7O
qkbhyYtIvv7xFgCTivY5earUZuBRE+cskuDgpw9zgyVeeSNfuIduGe8WbPJz15M2hkGPiwwn5fB2
9aIqOGD84rDmt5+rmZaV77l+tV6l/sIjdHkmaqZWGS751stTxleGbWsNFtgqWmCiI7MWn4lQBPlY
dfUCCOKbo0OJnjdiuaBlVPuoWNEXsMuaoPP2UG2MRyqoBJHR0tyrty01418Aa+NtV7gZXgtF1BpO
XJUD1TWggEh7jRFqG+lQajtbBHI1h9z3yZdRGAJjjOLFaN3IShMnnzFgi3O5yGoVMLfHnQsD2w1P
+jDkxP+L7lj9f7vGdgQOcA7WvhV/joh6LaRMyyPys2Km8S9/k84vd6NFxJ+NyolpfU8sA/XMNjbM
uhbLyuS3U57JzcWJtkXGFrgTFFXROFLNcJfOOYHGyKqld73egWvM0v99O5vSuQAxPyVRdntTJqV2
79FkDVuTcBidM80fihJqlmmoSFybqPXO0ZFgc1GU1586dRTqFF/m8dvQwIjZhWBDV67SvJB1V5mu
6aoSA1E6iGLQqHt5545OtPog8uiiyT9qoYQ8Cmfuqhbhebx8p5DNpcPsy8yftmOGTRC+jnOW30uk
Usu4oVcNsd9x451aCsYsKd/OTbr2YCq178LBfi3QYIgH3UeIlgokP/Wd1K99ORAtxmYD4YPp+dHo
PgwYdGtsKNCtCfGOqyjMjaa07mbxQu+lpAKDc7XN0/e8qquOmKC+sjnV+Duq4vwV6h8yxc2iRc3d
4AB0eMaLLBKIl5NoW8K+DeZo2gi5YCbz+bAkLQgvOmIR3LAJxPfiOcLvdAGxxhEvVrLM78X8sjnb
p1eq8hwNJ+laAr4uS+3XKftoIPipdLCkHVd/P9lci+ELPaL89migcFDwBqRlhVhqa2LLMBG94nns
gXPzrRrJg6gCkfduatRFHNw6DT0K8DVv4nSNhPWAS8Fk3LVwoQtJPKVvj15LzE2ZLot6Xmh2xHDw
8g2hY9LhmQvjrH7wCoE4aHpUjHwUPlVe9rK1GWmAcgORDF3ae4mbFTJUT4qkTx8cRJiIjrI4B2kC
V0PnjcJLy6YQZ2dHyv723id2SUiwfY56fCPt7omE0F0yLY/s+K3qnI8K4kRUo6d17Ca6r4QsdHe0
Mfa8EbP4vZuBpIcT8TXFmy/9AWwJwYz431IR+AXSwP7EY+KGQtovV8GekcTJ8IsXTIt9ykSPX/lG
xrAbAP9G4ULXw6i843shBwHVM8nEsj+kcJW39dy1lo2gRH/igtqdyCmJMUy6hbRPZoK+baP2OFth
xcA2FTJqWU0vM3luQziQNp3w0/fOOxb9X/Un65xDEN896qVw9dQicRHSLMvLAzM9VcLSvl+3RDXu
EWu5n923216MtoJiyGbICdv96g+UjzJZF7GONcnsgmI4CeulLgYyUqelfBVLugriCCcnyzi+ClOE
HPkQ7vkcLbys/MSbeH4SN7EwbvHzaesZzGv7nQ7QEw3p95hSqF3e58N8QEqRDuH1xv1e9Ru8sFj5
iIB/Y6Tm3qerNPPU5B9qSVVcK3YNYhQYEscMIlQlZl/FF2xbl6tUVB83Dv54wbO144rDYpJVZfDi
NgOxOje86fsrUuuqXreKrvtRe2M8ZbP6lSdDmBbp9UCb8KpagclKXUX77AN2RAaXOBjeq96G523Q
X7VeDUzc+Z9Eogv/4gAU7A332+IqsHhr0rrVnhkZv26Az/N0cQwoiUhleJG+VIcotXtMwvPIbCGS
nr1RuSQpENdfVsA8LK0675v4Ykt37QPQ6aiYOwtR1lN1gKLwRDbAHAnTEkD2qPsdhjUc1wgn4sn6
YiPnsp52Dt0Lzs1W4X0Xq+yFcVW3ySCv7PQPe5E9kx54M7Xd30SF1RRmM8fvmPyh/L+lV06ryo6O
KmSqMbrNWQcF3PPLk1HDfAnaswzwxylwuiq/xIWv+bAcXNuA3daatrPJJH7RCvokm7KfWaSYRjfs
/kdERXiMwRRZepTxks5blKhbYQ8AyxcnVhQsYS6qFjstjnlcLFxLY7RbIRiWty5qaGHIJz/U7QWL
6q0x+FkmEF/wq6LGXMGZ8eUACxeA+76PyxRAxvhLdjLmlXzAEeT0TDINtA1+jdMxyAmZSe+cwAqm
7y4lAFZJoiNbPyFn/NSN2+GxvBC9mSV/qjKOyr7bIABq8RMomQabDXkTTb1/9xEas6Tk4Pq4m1Dn
LQxegYzVdrehU54COKZuCFnzwGv0DHcKgBCtNUnp3WDipgD4La5sm/+xNpJdq4zDlpEmgiqXmeQy
J4pVdggqemDugyfSu9/jm2444hMx1++lIqNq+/XkuqURozdhQHbivTync1crb2VtGnVYOBgcgEHg
HgTLQJymSYJjQ0WEHam5TpPj76xtB2qPuGf9PxU90A5/2myOmZGCGBDBffKyhxIW9W/kPZ0qReza
J/zBGT1SV65ZVHbPzZqqWELvac+ekCA2sIUY5SaUGKJRASVRfigx8pP+wsmEtQ4waabnGTcYVLEL
M4wZPB19o2BXHo29JxDGwNKGRGBPgSSoZaVoe2EB6QPUOPYfU6q4X1HRXcyN5V9RzGwpnNRw5h3j
86PJhCIuKL7YXws+1AIvt+5cATwnhl3NnS9H89BafYUo0s0cy2zZgZatMh7+pqJnB3UbQPdXtGbq
sKSL6N76/1Aw8uq/gklyWDwZgvzU+Cer0DfUPMZ+F4ceTABBdPOM0PascF2S+V5R+klWQit0wuSh
c98jEZM3vUPlnn48dasWMSZwtfCjFw0ExQ6Dd81ewEjqRIApi+WzE0EuHEcM70hZhANHTOhPlvMZ
8qfMVaOCeK44s6WfleqcZSiVNgs7TNx56HwwDx/izsA6gqd+hwO9rbuUqUDZmKDgbZi8vt/C5w6p
zMECn1/Xx6IlLz2bxLvRx6Rxz5DlndUTS/fS9HZsDMfsXqHf08uoqOdP1kNN/nIaE6F1GsE/B7U7
VeHlAbtt05BZLqGeRt7cNmBQbam/Unj/orUxyHDpaAmx+S6sQoolgAhov+211ckUOSnvHfypaLlQ
qbTugpiaPCULwvH0zsOvyIDziedNRrF+cfswDDlVrXPT+xzjzOuLGn4CnLMz35HffX301HVavJtr
UWP9DDzqGWTI8erYeeHc6qxGVVkUUGIK987FZoaS11h79HCSj4i6CGDmtwMKazZOmSlIUPW2IHp6
evM1yE23psbANp1YXbeMkp8KXeRkduX033O9pYdY58TqduryxBFCNJdSioy5hdrvrFzVbPubXtTR
q58XZN71tn0N5a8Nij7i4RoVcEoAz06AucYq2wWgQZZ8a4Ru+eRATY6BRNDinK2UyGUqNHAYkZMl
122DIWO5wePhKGuVWbixn7mAs4dA5F3nFYP1XNL2UZvyYQfT3Xzf/VNw8nqffbNx54kpOxKSSnDD
xvuyMnbTSLJNAM0NqpkwZPbaJBMJih9FQ++rvJKjz7dXBHqTctkyqgTlqmq6Ujp1JwmmUojFijV1
z6ROa45rx883ypJsj85S268ycWzkUmnbhOo7DonSzwKCg53aoRq6raiBL1IdawuRLNl3tckjZbPt
QFtDhk1xm7MUtGCR0Cvhtu1QlfvyGNz/zM3gtL0bcQuWKkWW5s9MOMQuE2j7vkpngdlqr0yDdJuZ
8rrqvAGTQP251iwoN3JDfcPREEbO8Wt2QG+xdwVrKKGBBROvCUuhBuLSzbxNyaNcPggqKxgk6w2O
Teosp/qiLwWgn/Iq4VpnYceoKGzwAX+u4TSc9xZCdjiBcayZC5kUWkm97mEJ5tqPD4yoafK7sS3A
MImfGwKelYEHwU0g4drTgqfmELGEGIJih6NWLnMcBdi7iD+DpFKxUvSBpFNghLjkUtGzw2OhPVxC
3Bo2vf+cpqnXmEddjbn8T6P7aQr/J8nXoyTNQs85DaSxaoupNi6XNfVskbWVyYdkDx9HVlkzlO5P
+7TCO62MLf8wMMyuqrrpLC8I19agWPV2Ke8wQtY21XFpJok5DGE1aA2kj3FqSDW5OoMw9lDHxlNd
tyKBweLINuB9oRkXv1kc21Csn4XYWbNG+nBnGuzD0OJxTg7LnWFKgr6bVweTLvNO33nj3HMtKib4
OkjnNc4vNp0LgU4w14xuNZKP328lWVhiEKdiBLbXhocSKyI8/RikZspTYKCLwA2DlvIwbRRIyeu6
lGhBZTqKNBkChKcs3ljcC9UBsFPAJk0RkYZdLUuLoEhEvVgKFjriRte5bih2S+By0FBMeI5QuybI
w9YKVqxH+pyuph7uPMqrkWMOA6dBVhlOJMvbVoPf8MekIKdibOY0RwpVOD8YKzqfOyPs1NC3Jk4P
10H7IHDD/3LH02d+VKl5eeCnx2g5lLUKruEOmS64eZ1whuW24TrKjD6eNOnT918W/v3YhzpqA17x
ed7j+lUdklNcI5tZX/piPIS0Sqc86lR51dWSLwIyMaes4E32F778XT2SNbu5vXMtEg1tO+az5fi3
JMjuxYwL9z+NUc5uUC+5Lq+6QE9VDpAtA0ptx03Dru209NJdSXqZ/dHwAuMk9HHywRdhuA8EpOQL
9IFuRnV1ZzNsOE8hM27gpqvRwwjSgyhka7Md4X2nkyayC2QqAflNRDPkF2Q6Q/t7xK0w/RhJxbZ3
5+cIvOqu4S5+J81ZVKtoEDmCCsKyQR0WboOp9levIB7+tfocO75eyxP/RwKMt/cFq4D4EOK4o5Qd
O97KHuzUW8/5BR5cYZdEviqhN/mMxZ4VK46r0wRbZ+raYD/AQY7c/NoHh7lAdP8IOFfnU8Bf3uPg
aa5ps7O0eENjBdls+FTTvSUyONTNMbsOffXDcuoLUldJt8o8trqKsz2b2Lfu/1JOCbsB6ZJ2uCnt
FPGyuIBjq0fgsMTQpchb1IZZfv1y5ejlmFI/Iy/GEStQW1bJ3ogBWpxi4miLHz3k6qfAapOtApAH
0TQcYsQ2OtEVufR5VBMSE2OIKC2jUKOmkilkWr1Ovc3NWhSSiF8rUfYLW0/D0HhgQuY4Qy3mIs18
JvwYgTBtkFX1bUlDJhQYQ2BBI3Nyxg4JSzMwLVAlpeE0VRXNlfKlzt929UDCW9F0pa4AEOH+BMfp
eRnxS6QWiAxPOUdgj51KzriskgT7DE9Pkq7FetGRLezwkz26JCO5GCXAlAokr/fb6OQtEkV83n+j
UXNqcGKFD8KqR+8f7ZkqpnnrQtrn4FM/Rh8jOXg8aFxqql+bkP6PZBmEofioNIV2sns2zvZWFXEZ
NeDl4WdqbGmzwiglXDwdGQBsLAWrdSGS+mwVz/dAf2yQM7xvKfWsSnLb5lggLobAEROdIrL/nRcH
Ki15I5VSsGYSdzTz872dJwtEhC6rZ2Vzbqtbn0LG87McrwMhs7rGlGdheGNCMdX/AXkbcD2G79VJ
Uyw6QD/CnsXGP4tCLLA0L6ePSu5Ca7erQEXVnOOofJSxWdvspTPMCRZdPILH5Okw/Qbhi5eA+yCC
4J2/AlFuqWSZbc1IaL3pKKcB8V4sd/m9DLkp6LIS5K4OsGQCiqC4Z5WJ2KDYez1b2O2o35VuYvzj
L7eRVXJHbZrq2K7J+kT48QDDxeEEyqfNN/Zgitpq7D4HI6Gp2FmZobmpkPRGw3UPvE5SQwz8BQIx
vV/vj6BPDPCwqFg0OZo2ZYzeQNN+UZz1O4VsuqXn8kBW6rQDwywB+u6TvztC7fEkKbvkltdGJeMC
E/FUx4VR+aGp36tyhW2X9vJH+zYdd1yBPHuaUoH+A+90Q60roStZdpsrRGk6INA0hVAWQGVxjqt+
H6hYmvt+jTCv7YOwBR3WvRrRyRKSDRiOU9VdXeXkhQqxMRaKUu9De7HYsIJmXK4+34uQ3fZDe8FS
3S7LHURxo5FB0vQfN6FO/tEaKvz3cI80So8/Nb3Zi7zTrNGa0Wonvy6nLm7PF8ERtii58k/imc3y
gpgMHC2vfNZ9PY89WY90gV4hMQM8srtf2UUIBWAYfuhEOc7HYrNWiHEdVeZwr5ysumIqibw+NRe5
/gJsRb4/UiD1yhMgPKJV8MjFUE5uVkiUYk8F0odU7ijqjLxXRfI7Rys0nglWCzWPNxlhghZJroyF
wXyvjU298SSyAKm5Kd3uS4fslTqLGHO/PAOFqwvq5cTJfji81/SIP5hz8PikZ+/5sAoMOJUbmNdn
0AkcQLEc0dk79bA5eLUUyDugmZ4MZRfep8xc9aId67bi9apStDMkY/x2Ac/0EiVti4aJ/kNYLalS
yyaLMWEN+Ov2txXLVBEkDf2I/CX4lBDeOzidOTD3uLhLfURyCIiNPn9vlDyWVUDOTYvEHx3MreoU
K3P8jYVVvTilUO1mv/qQYNBJoH8CDMSLPevnd6nrCAciOPZcWeD3AnoV2XWOkp23RKdp7Xi2x9Et
r/hwJO3p6PJClIKI4WF9MXHuFc/VKNAD11SUCtrFjNWMyt3widDyldCIvtnL0TOL84agoPO/h6Qf
tB31jiNCecO5V+lMCq0XhWZghSp+La5q1ambAYJ/C+w/P6eeEeWrRiaSZ3P+0RR9Qa7ZlEHbb3tW
w8HXt10G+vItNbBOjNEgok/sYBCINhNAF9sU1pvMLLyMZYzXoP4+ccYd84tHWeifZeX8lO5lpdKu
s2dYuxiDepBUQKtA0y5qwcVBYH/VyqmcpbsPVHv+hEzFzT385z8KjEkX8pv9bJc4iVDevyaB/lO2
h/PL0TUsAF5cmVUCvSFCktQdeMcIZ4GolqzUIGrNd79yGppWbLPYNP/FbSpa82R76OfEnYLVBKsl
6huU5w8LDbDtVGE+tSj1jIAzAbcqft91AsyPbqREb1c1yX6EkOeutlM59p7UlNl2rzX93Us0/d6C
KWgPusjhDSR+m4jve5T4bkJsL7Rni9hxd6pUCtDsKBOItKdxU+n/OauxzvZpw2D6I0QZqlpIwfJY
snUH642C5DEEOFLZ9wO7MaifFSD6/9O42tvjCItuhilOl7TkdynnzP1kAMZLmfeGxZhJG0CVGVRL
RuL0i3zxzSJ+1ZwSszuywIGEGOaKdADQdbNmyR0sr8xU7QY6FDYtlReU0Y64mFTy/9oaDe7Brr5u
LJhay+F91+01AXUw/ZyPo93iVFMdUY0ZEq6ETxN52dyvXBdA6J5DPw6X6j/tK7Xs6Ec1Bjdiqx30
qd7kY7ptdjcgikF3ZunEIlOAxP/GEX6lGpPU8xr0eoKrU8SP232Cbih1aqbgmmSuf0weaPKYa+Xm
KykocmnkYEAV6kuWMEAeZp8/pVV3DEnuVwZLFva4zdvt31Zw+KiCIvcuKhAVSgcMfK3GpsV57lTv
d5oEN5Pv/YrnpyULLk/hthVh5wShFNNS7VZSzXwVYpvt0XyWSBqP1z2GYr77PzjBT7pBKHPXIbC/
JBtMR/GARd8o+gb6Y/XhlRyCsAJ2ZKsHx0YpUw6j133/dhwrOmeegq125MP1R5oFYw5RfJmawjTx
rcC5p/SvDYs2eFyoO3uAvO6SfmFZ99GTRb+MRR59t8V+o8MLq8Reihf2WxVwdTSCTyD9s+ysphMP
BAwkAaZxUOJrKVqkOdlwI54m1d844FE5h1m0uBIDwGKdMMGuvH69v9GsVYV8ZTcwrHL0WGrWPTEd
DDmR/I4JuMGZLCyV9tq0iWRonLPabMB4snU+KErdA74vNUULHddb7syTzM1xlFlc13dcpcrcYQWl
cVajVieHUvtLWANRtPcoDIDGfxBQAeYXkJEX+5VB8RPuTOqU8tNC1citKr+QRbblHYt8fOMN7eUb
oKpFCWCiCy9R2yy3ToYL1o/Mif5u4qolmWce+5eemXl4bRv7mi+SCIdxTEHU5guf/8FwK7hAnKSz
RvD9J2kxkoHj4ZjCvRGxaBsRkwrJDQTmkkSp7bD/yqULEWRo+fxtRs2GIeIhgJo85AcEavUBMyAn
GVL07BkQRDzWC2LOi02uK0CmOzI4v64WGkTCBPCjJ7RuvfFOfxCL01pd8qyRrhuVa60cHy1xO8V2
eaatBAcgBvPN4vlDYQkeUswIK4xSm1Ww1zf29qffjMQX5I0RFxxuAiEKDk1wU07tf9eOFJ6bBVFC
0WkDxonlPQk11HqDkZS6u0hPhFGP7RRMTE2dWZxz/IVbW/t+6bn7h0Lf9UCy8DqwrwvlIT2AujWa
Xv5Fb4vpvsMAa+wODNa/KLjuPcMzCpChuwu8kJsai90UJPjSJEYjmphv0yOHV12IcJFkiWkQ+RNa
dOdGb/eVeQHMRj271QDYw6oo3iIJ2jANNQb2Tq8N4FPawu8r5G/E2zCCooUfE/WvNqsRRiIMvFqO
AFvxaweJWW3MM8cLSUiUrojysTR/2GbiyZNd586N4ZoSGVxLk4Nsi5RF6C2o+EJ0gGTwnFbOwqor
Hcfdn1yNsIgxxUFlTwWuJ7jYxLRt9mjznZHn/BoK8UGxqQLF1+3jsU6CY+UQosmYgbOKgKSZppzz
9dpPl7k0rJDuSxOmgvUzAwFxBFqJtfxZgTkrwcDJgf7D5+zJ9M77KL/te8/yarA9gMAg9mHt/kA7
L85sS+8+kFDdsB2jOMWTvuAxqDo/XHmmjcLrMYiim5haQyGYmHpDHiXdQhkEDOQBFcedx3BrWbtL
I+5OQjTffKTa2y7rnZtamNpqFT7xNZiNrLAd4bw/QSejqKlPmPeil0cmwhqaCPQ2nAQ+b18ORrG8
kcg85fVE807rlExKrQzQOw8PBBdU7Ty4fWgW/cU5GCd/z3fSSqANl74+3ZL/96tCiGmUejlm12bn
qjY/7cOkZaJDiE7g4b5cFL7Nb60qiwtNTMPI8/cEWif5iHh8aJh+t30DWZIHR6mlasqaKyXNO6al
tytB6lWJSRZze9knUW9WccSqtE2pVnLrTnT4XcMBIbiDCPoDUfN4UE6g09sy/ouag52hj/uO1Ax8
I9XSF1KitJ+erMtfXuOitk1zSrh9GPeWIgA1OlRp+sif1IRu3apNkSTZitErEduPOeoUc17PjoWv
Lc+LuWIQnTaHJpxMPUNcbrpQSRxeoW9HFwzxrCUJFa2sPmO5Z6t6t5jqGQoIAw0qW3TvXu71QEFY
Qdrw8/K/GBvOy9eklZk1gfLgJCd0eoZ25BApenrhj3kS/EUpOT7vyzPYB5u+bZEgoG3FQR1L5fjh
4TasSsAawByU5r8VNQ5OGyY2nfT6Zwji26YRLke/2tGjWHwTmLVz91xn0TaEPSs6o8ul28ZrKLgO
Ds+PjciSdK2lONRCI+Z5D1x1c95yrtJWKsZ2w8mWofsreXuDvGez7ocXixZQ3YzQPzTJ1rMlKPs/
3kWKN6YtC5jBYWGDzlRhXyb5+b7c927kULhqYkpyZJa/6l5NAiswxsyfw/mWNUZ4PfK2SaE7mQ7t
7MXdc7oJeUlDpwnCnAe2Kbz9QqfxxA+Z9nXRVZZ4jKur2f7P29rOcx1MfUG3p2ChxpXcZS9tKnx+
ZEdySGN+i5eQ2ygC7PnPWTjchON8kvRbeeSYJZUY/SvCXnDcqtlVefNk6cocWPGVGd6T2JaL0TaW
fAFfAdQi34zGeWBIkef7wct3IHQ0AE0HiF2Q656b3L1A1ZZ5fpMA4D3sXNw7gxunMow0dRL07+Jq
1HD86kMGTkQ0XV99rsjZNIgZA0ZUmte74vOPjV3UPPOhZKI3rd6DYiF/uSWxlXblE9ppbYPDNoJo
GXYU8Ai/e24bYNre+KoFIw5gF2ysgrGCEfi1fAYvGCC8Hr6vtgixf5tPCCGi2sOPGArUwHZvtP22
P4RAwkBY10SQ+iKNCIWKn0Kcv9/gb3QunSHJebnrHFd06QW7aKgJTp9vS2bB0ryosWsUPEATYuv6
EKu76EDAIKhc1IWsyyxmf5fsSfKmF2S0Kx+AGrKtgbXHdw6cgmjd7IlX55cXSAnVjmq4Ajm1JyTJ
EdAAV9jQOQTDU49mLV7jBfaBjiuDHTmwWbRwSVXi/p0O97aPycs5a0CHW7QU7+LJf8ayPt86sY6A
klkNAVDObjniBmrI7WrkI/BAUCKpTmWKFLjnXdXEYJnisPNnzXBUSGN9GhunOUKBHB7olHfC2w6p
F55Zk49A9F08gblLz7o8s/KCu7ITwsy8gW63evIJBx45FL+NCh5v+pE690QBVf4BQmlGhVS7MI9Y
67hv6Kit52VHqx0gdTxqMEVDo873UBwsz25g72jOdBgjge08KSrE7AKOsbWX4ciL0P8Ts1sJdFbG
x0jUhchexIdIj2oagCEK3g5K6v1z4iIknNlKQIkCxvpx8lJ3ghaf8lF3dgK+C2ALKq8hBskM2FT/
yEl/+8W6HJrJKBogNIScNbSKOSU6sQLykipkSQlIUIFTFzwuX/dLDMJe2iaGdwtGVSC19rSATLhL
6OWX+YR8kyC8qG9lC9mNcOwSLOSRGalusZi0f2fTkAnEauxFa7VP5UoTfpWfD18vJYwsG/kNRG95
m1gMf9lRG1C3Qc11bEGOewQD3D6Otz/HR3l5Eq4upoAX3FY2LwOw+iu4L83DiA4jj5TUDR43EQf4
qFJsR1tNkv/9zjZEBnjw+BNUeYiCTTDi+66Ua7sNJVDlerBigfuxFDioeoXOOdMcer1f0SVGYLiJ
v38GkcAhLO60lwpw+conYNCXtICq2sr+pmKDnbfF/HGV4GlM+Ys68Cw1ZHTpmBqx6Q0QUJNpXDOQ
mFPh1pkXHbMYyQIlGjoMTPuX2DUkZaXWb4d/mzlw1to9VxGYM9ud0TKkXn8vq0HxX2QhMrTrTcRM
9H+3/bb1VA2pMOL0zm6mKWhpgJQTAHgQxB0OzYDBli6HSpoogfp0SSxmeUoMLbBPm8ghRswLIggQ
nfE9DUu6tE8k9t5hbuUb3sAMbvwzsFXsmaalHp7yxcsQyDOQP3TpGYVw1xA8VJJM03O7au8Iez15
a2cw/x+NG9cSTYQLfafgkjchspSV2ldacG3sCjMd2gs5yIaNcW6IyTOF24RvVcMuy9ab/YcogOV/
hQq/yQxSLnwFF+q1y6SLoiK6GGyAORisgH0AU++hWY4haIMtd/amYFWb/ewY+JXdc4tcNRdmslIn
+0XnlIJzERrMEjcoLShqRMTMN626LLLE4ZSPMVF7/WBWws9aylXKeALbJ3MQQwjSu9ScHTLHm5DG
d13hnlUPmB215KA+0YLlP/HuEY3qGMmT29QSDRF7qui2aUAkt8ctgxGzLHX6d6IF0Vc/lqZZH9tC
TUdBf2IIHbhvVrqU7DyRelWDDPNWSeYDOz/byujZpxHR8RWOLKBouEh/RoAxribjAkQBKIxGb67x
WB0Yn5K4U1E0aDYzbN26Ui6FSfypUMktbyBhFGypP8S8ViDLWFvOBEZSfWCNz4shPSzV+4tqnKti
b0/nOAC4fa5kiHCrx/9PBbi6wtyVCvTWOk0DGjlCHN1R4ah0eSDwf3SNjALpIGhJeL+3DmnnYiYP
tlFFlb/+2Fmy0bMyz5SrxmU0Hwd1qLCU6a9tvT+gzwt30klUfSdqM4oVJqzPRbRPDApafymQP/Fb
J7GhVOD2ClSb4RfMMHeDJgr1YbhOeNpCJckcVsTldRg8pek0ULdDmEY4ppffwlre7aI6vz8Puy4e
BxPOYfg4C9nHYoAqN2MXOHe+xgi4tgR4go3aFTfehFD0NgBXmgNLyRtMhDktHUXaoE8E9hPC1nev
B19BMa3INof3greG3HsZo589l1O4ocDLToSXumXh9oMOUfDLWuYCVD6ygJI52PzXFLcxa4ug7zef
1xnkabYBTa7nFgNGBbE8qM+A3oBvuOz5QBmXfbNMHC6dojozDM6J6DwiCr3LA37I9/LT0C9nXzmE
DLt0UhrRgeai9paqGyh/TB38OizgNubHjt2uTdjWp7WZc1wsxGhOf40zeVHUz+ol+EBfecHdn9PQ
6EY6XDFsgycu1DDqdJNuPwa+VXoaqcZubzyfd6FwXrnhLCPku64LjoyQHyxrydgo9dn+1qqdOSB8
hBrGMAtwUhDxX1LZY42U/v1vBEb0bINX+qx/F52N1BjEAdmbJN1IHunXvMiIp+p36vg+PcQWCpeB
5c/5Jj4/p5m8zHQhNdw3oCT2YKqEpKo+uqCWM0tQ7IXQ+3OLJ4VLwQb8kMzF3ehK4/jpwqRd+cjC
k/+0ycCOaSJBN2IxiVi/fXob3tAT9NkpYoibFbgLXoQitrXXr1znRsX1O/Sr/i+6BdSF5unwxm1Y
Kh+muMALjMc2YRoZYeZZN2zBESMF776YHkCYWTXxqgs+K6ExSIFsdp7aMruWY/62TXhexoUQE7Pl
9MxIqxpYpobXoyqIwHHwE552dfCNPk1p9q+sfV3yZgm4UGexU0wo8/B5BLAvL++raU2Z240ys8rG
ggPyJqtdOSt2gs7NKCCmCFNAq9pd31rLhC0ErdUzi2fZsEt7+QKolZRBBxc6cWudpDxVVLiWcQNc
QVhxonnF9FD92aO1mNZFnqoVta1zJ7XCehlqhnfoNcXjsdcot98JC55OBglATQmr+zpnvChu4CRl
79W5z1AHf+RWFcUplkzaQDELpPYhxWxbJidQMIuA4lbOdEz6dwKUa5p7YrmVg43oqwsTc0cU7leD
QxSoqDYvL1cwNo5OFjBQU/hBRoSottYxS7Yqss9OV+nc5qw2pspjXkIq6TzHopRfbxtTi0iB6r1I
JF/HW77vGzjocDEONOsBD9qPiMB9+Btkv//+ljU3LfRr39uFxNMy80wwmfdb87C9r9pEdVjq/lkF
rR8/d4CwBeefYwbKGjXLvMIxh0muqH9ev2IW+6AAtuSedXBxBGlSGCv7p69HD5m5/DtpJdWv14SW
nu6ytNSap6oB2qD6xEEer/ZBfuD2QrYRDPDsiIqKsA8z6sI2JdRTILyctHRvP90F9EhjsI4B/NEO
bpymCgrk/xeJFiIxI2p2XtTdKJYW/S7InwyNBUmcezVVJLU5XCxeMH53ib1mOryeJQ8cd5uRLlMj
pSB9oCmeCT5cvqIny8Sj4sf8dLAciux41jsMqXQrZEZYjaU9LmUOKkOfOfigLPKn2BDppTRv0ByT
+yAauv7l7nCDInlv2QC0BuWnhKqPbWnhGKNeMsHY2c8PRVRF/67n4tCso/v+RpSiF2kZZYBahLMV
oXeKwNXEldvbjYzDVFVSBuZiIZ7XIia00ryKMOqaKDujTPB9hu4Ba2rgM4iZfhAshmaMjyJDSdR+
PFqqt8keHC5WJC7+dhY/DeYFHNPgjt9t2HnIa3CFOVLvhugaTlSKjRMZ+eeeTCaXIRZy4zGCTI/K
G/BE1kb4IzR4hR1cuGc855sgK2EiTw0P880CrdbMaOEAr17gCgFr5LBZ48pkZPKa/WAsTdoe5eNj
tStpyh5NInQuAheiUyx+h4OcsEDVsrpVD3h+xEBH9kAY9gy9LOe4jQIWK9t7s/Zslhhsmm1ZIu1x
fhf0+GyxObzzbMfwbo0TZY3Xgv8ZAPV3fywRrHlJ5SEhQbz5LuVpymMZsqV9Ox2/ummqk0pP4phC
cBnaEVTaxg9L7MBHuqpBeoat0UHxZ6MdaCSoQdZSYVSnKRzaw6VNBav/nN2yTnqbmQ1cPrQcP8cS
fl+9gYILmfIH4kWO4wl9WNUiMDgLnOZc93HeIeHDK2aDk6rOLNhq2p5WNdBnjId1jmHdup+wu92H
o3iIQzNuBdsrWMVL/mc7bZFYgMkqtaI2O1t+rwi0zrBIgEcDqQXSLtcpFnkl6c5Y80hH+ggH7/Hd
N/F+RgbvvTM5xKePb3prAneSEnVVbKr7k7Wo3+ll3ulcoS00276vVodHpJFPIlT+FKNv29xuT6bn
IaMTps/TaDwDmtDFDQcmel+3idb4uxq4cEqu/APQGG0RQIHU4ejO5Zi7qgZZKjyuVN9LmYydE8C/
QabAIF8i1uE+MqumE8F5rnhiWIOT2C4IvY9D+lJrcq5STsa9T2RFlldcu8zkasQOpov2QHRZihuR
AK3ZzwQ6pU1Z7ESJLuRqt880u3PuQzMDijoe0ujIF7WQAFkkY4YzO+yzReugsmXriGmhqSdckezX
QU5A5Funq7SAfFZYee954kKTK60ydYxuL74dcKgg02WlVVvFjKaOkazqqpKCTNn/Db/G+ISIPuta
HyHagGzmzAXsGIdrX0fhSL7EFXSy0RhCNmfCdkt6L3h0fXa6cXaYDU2AmKjlTcSRLKWJXV1wGLTO
DknPsmJyH3co4oiEhtQ61kmD4lLky04Ewid1K03ZForR0rSXJiPJUUh+T4P6z8fQ6/P61WRsP08I
vj/gjPSsuChTW+V2Ctx8bbNHLkYB+hQebT4CI4M+K3ZZDc61d59sKzIfgIOYnbn8QYR9vDc4w2LW
RgTy+DRxWCCXiChIZqPihD0b5hJRbxqUWYuSEJ+PUqqhCBbK/d1XzDyCgFa7gyMXF2Ii+6vaZ2KV
Nl7ujWjArAcCTirDTM0L1WUQpbxECHIqPxhJtWbjDHEMmHoZd7cr2lbzWZdrV7yn2n0Sl22OJZLi
sOSxfUNtMjtqPEvBF473i5tMeT9ezyKhDp6pvxA0+IKhFuv6CvhAiF+G5H9Ej4lFPKSLZUpPeAxh
x184bysKApBA5dDMvhW5M/CRgCB/Xc9PLxc38GyO47jJMrHKRZkqtj/VnjRGw9iUzTZZeJ2QJh1k
BAa4FiI8Hqq4LpfjhhfCQd9W7o9qdBVNMH+Hu4sYofsKBIx4/+SaE1kCCiaEU4gvHZenYGFGeJNo
4oTpk+oPPEf1rW2eywLIHg9w2hh/Ubj3EQjoLptiW6mf506eZoHNLD8AxYe5BSDaFI0dEUxUjwk3
5OtTPQwUKR091ZjGMZQMFwVMmkkKD0Vm1c+oPLZuU9Fv10EmLSDjxnyCZe3GMIxjrXNdGyrkPY9f
5sFuDzeEJo6Wftsfn8+9yScmZg7jlQmocRyt/YkRNVUZ2c+MSmk93bjKxZhL7LKq/MjwReLJ2A79
EdrCmPL8byF27BF5zuy/IerJ/vU5YpT1MpADaCxt5lp03opKeOuthzVJKAPcKOtIG0hy0SVM3A6G
9ji0C5I6VwPYWDGHRSr3UE/zsc6aSiGVipvfpbzZUsd0EQDNAmXIF+cve27mpdLG3mcFYmvdLhrF
P9QPqBBoVgFCXXRkIoIk9YQeXvLjQBWNYCt7cZJ5G1emS94j7l4LnC0tkW3UxyAp1c0jyZ41kSgn
rz0J3QO3sWFFUdk7555UGeLNCjbYxUOnNtpUEresmwKYmJhTHrBk0rlrvqV2I1KYSiMiUFSV2CrX
8BsiWsNxf6OgA+WiHkvoMFmR4nIX2Q0W0Oy+IcO5RxINdokOEQcxcOIAlybmZ/qsfjOzB2mSY5ZY
fctAW+QT0NmVxG4WjOtjsTlOrtBwBsDkVx8kpT8/uQOHHqJNFDrpqmVPAAHeUmAcu31ehWTawe7w
uiopDh1TLTuRfmxAdNVyo0dVWlhfj/gFtNI0inFfe/0uLLZqQ1oKaDJM2OjWtegpBZemvcuiXgHi
JVTqBeGcsGQlS/ISi0GOrN0SxJ00SZxvHEfYr0tzSH6/uI06esDX3Unmj341PwMT6XPWi3YGVPoI
uz8J7Jpxyn5yp+nE4BodVPNOBlyeOq7DU23QQLUY2gXpG3aEzJt1zsfUUttGkqlLPuBjyBCw8eky
8bgv4+9uV8bVeO6TLjW3PMi8BV/YNCainFte+XmvsVXJ/yygoG00pPOYcCynn8Xb51cINRqceQJh
S5jQernyBHqmP7iPGRQiJZHdMAfYv/TUEGzvjI9N52p1d+sZloaaji/tCpkgKQI7bDCZK72SBw6u
v5k/CplkXzZNG3s1k9iBaMVYI3mu2qxVAi3fgvcu53Xe8cbjHJUl5EJIl3YiRvyvAeOGR88PK9Vi
75B/ufTBePep1WUk+tW5ZcLbkTROGpJAecfB82CH8tfdacPe7zZJdUFq2Ljx4Bid80ne6l9Nt0eG
y2AZJi8C6hv7lFB0TCA/MC9F0JJET36wy0y9Y+bZoD6vfOmCyESegaml/StnEFLOSnshJR2T6o6g
fDoa54FrSr/dwQLgn1Ll8fwJMhwHdsiCCG5c3c/iAXL7I2/WhizgKL9HMeM2zoOsGspCGiSCC7vu
HwKmnK9j6f9CtgjeVcWN4TUkJgKcIvZ2ZX/5zIn0H5kdKyX4/KqbWod5UunBG498MkOhvEtgbx4S
6w7kPnf+wi1i0C9l6UxXMcN4z8lZwR6FFh2jM0hThn5M5mgy1KU6vxkoNfZGmWKVDL6z/yzri8p0
yOkdXIy3tWadQOfc4HJlobQasAFIsbopRE2VwuPWjxWCZvZhVy9bTh5qGStn+ywViyDMxWBuE4Av
l71pDVoGSBc6WBix1J5sPfjFqhlVk/JyScFQYzf+Lk2N/jCE2jC7VCpnmGVGrOsro5csyFKgeD0Z
XPZFH2HKE6w5d3i4mboNfQyYSxOFI2B6xEvkhL0L0rVJaUBOQQkTBHYj59rR+lTsrWk2ycg6ekQ+
GAknNLQmwFr3aQJE7RINwgf5e0k5OG2sNrEknPQOSiX7UQJ5PvN9/9wvLR+YVuSoxQ9OlvajxSEy
jztC/wWDBSGSnw6A7p4fFo1z4mENg7nsqLMIBsO+mp2+z8DVykS8DNC/EiJv75bs0BKPu/6D+pvK
JXbYqirvdDQRJpZuG3Vzr9t1M9oEFYWMjvPr/LTuqk54SzOXFwEIQqprKNsPAS/KilOMsdVIX28b
3cIy1kwu7vfYurXShwAp5roEfxzoRTeVCtjGGFOvL6uhNPhMidIT8UrPsEKcNfA48oAuuhaFh9Fx
A6gE8hTrQ/VJQxjF/CjZEpIF1F4roj4HIOXjgs8ZFytdYqHuJR8hVoAhSPkDWH+IzZ6ARrH4YSrF
regP6ab82B9Igl9DL6VBaZZIQOczYI6OmtJx2WRERJ1888L5WpAuT9CMH8+iX1IbpVLYvUNxxHnc
2Dh8Ve26r7D7mXN2mV6ed2FFjJxj/b/4viz32waUnNDo6SsE/kA/ejKEEdvAyrSEOpwQQw67fkZi
RFzW3M9ELvHUPb0ZNxL7RuFxdx7/QHuI20LP8ztOeSmoMF2rq9qJNGPwZoD7TBNeP+5EKh+nLnBo
zeEcWDRcUKpvg1gJRkBm+mqyWFJmVpxcW72pY1TwIw2gTimA1aAEdkn5ub3FPi2z5caXS8iFGYXk
iBXA1u9KVeJt0HrsHj7v4v3GP/KTukQF681xVfLtwDgc7Ume5cxVtcc9YhO+DNQF3h8iwyehMw8C
xdW8cyqZi6gjMiubVdO6Wnj7RNEt5jtpIwOD0B35WXSEzPUrQ5t+blDDXhoV3KWGqhThZ5RGWjAz
Hk2u2AjTg8a4/bwZX3kLU7De8QFK7IkO6cPoVRhDggTwNmEswb4WpVThbKY4DmXfHuZUyTHuRKhI
xa3uzLEceOA+0EQdPcnFbJeZ+M1dXxru+bDUfzWhP7S/nwoXhe80FHj5NZugyiUd53fr4rUbvBad
y64VFELJicHmIim1ws6v1EjN7Lf5AZaZvPOM14qFn1ZTYbcsm9olodj1DBrhuz3yZkd+sfCC3qmp
XOuhU83fgJ9XBZxNQbu34AmFlVHyJiVrI7tOs3q0eSaZA1bLq4WQpTvZp88bA4YL6lSa3A0DMULl
0QcQdEd0QJ33/IFmKnMWXo0HiPqGRlnbS2LImK48MlV+C9YQzVwJCfqpE3oVnrFvkhhOY5n38RBg
pngpj7x21myrDnVY0uWC1rHVB2mM2c5jLBHfaE0ubgFXcKcxnb94OaoZNKNXr62d0LmUH6kiWLGG
rx8/lgi+N9NtdGLKEH+CgdoMbWJ5OEDnVA4jHdik+onUbFEWTInhV1u39KafTufcgxvvT35GkTQF
xo2o9R5zYkKgSxcpkZx5HqCcJAXFg3WxyW7sHVHpPlFtqCpx68U1k7lkJbUzc2OiDYIo/hLlSK5F
ZACGXY0op10rChkSNtMkOF8EwIFMn3YR/Yty1cNHZuZtE0Yps6XvezObt7qPtXsbgxBRWz/Ggedl
4DGSbDfQMHgOx1th7KLEKHCYCUq2Z3qH0oqR3+cFGB2rvAhRJ9+Q9ZsnYyj0yyjHjD9c2SflahBt
2vvYNx06YagreA1yyajLMRT0k6bZ6znPuCjAhDv5M7DYcS+WMypYhM4FsY7OuK4k3jXm5MH6vPIR
lkRec7GKTMzjzhc85+hMr+nyoITFWGE2n+JavrKf7spUvgFBChrJ8jQ0uqc8J9SkoAKEo4ul1yhX
lzpYEZLLQ/qQQBPW5KncXShzUcPr0Y9RO0qAo0i3Vkm/UjLpoHvImozymySplha9mbqUFj8gbLgK
GY4jRCE8UEPwM+jYoQtKNs5sMkLHzW8w4S+q0MgYfzWRJIPqpj8Zc5FscgFZSC+25mI5ukAccxIi
5cNKWd+tHw1XbHhrkaYbXDo7kdYljW5LEDN4KXZpVn8ZGw9s6CQPTuHUeI6CUYqgvWKoshIZUu1H
6S1KdviUsoOacHrKWe47dwI+53HNAA1jLlKVjqS8PE38cVGYwRs0ijTqgsWAN2m6pbrRa03/AzCV
YZx3NRDTR19uS+VbqTAIRwQ8IWMoqvu4D642F1/2T2MR4HMnTPCyV1K7UW9Lzpjb0ICpymppogYf
4GlLQe1KEA+UToQgicwjmnZ3zsw7/1iMnJoGVCEjHnjN7Y2N1nzU8LtWyr4x7lY2azTjtCnrTPkv
fq1OJG3FwDCdSjM8jSz8a3nT3n+vQIIsmQXtq3/VG/CkTsnPhtlhsH7zavfHCTYmytJEdizpkRUd
lmp2PhOA6cQXbwXiavR+Ovg24KUbvtECagDNvOvnvZGtslSTvpuBqZ2Jy4E5+LiVScJ/ZERuTvl9
S7z+CaBBoiz9CCDq2ElMdrOwSL/U9106/1FFrcB2PuB3ZEu6CGtRZoqpvnXP+h48U28az/gA6wqn
cawW4fkT3P6++6ndXrD5KPA4IA04ioQDlP6vwwMED/0moW3xNWIjtxD3F4rYh8a+JV40Xi3bzlua
QH/4Kx4Sc5SqTN83gO3h6pU5luqjRbQluzTHwWTJ/2K4tMSSMOvk0sh1K4MBpufooX7Hb0A3dV3q
UanQRMdA10LX2RITq2R+1oZ/kWeE11YPbiMZ7caiGlw3N0vD7QdnN9hxYD0C6yhBfw4YgWIo56H5
QiKQRVNr4UTKbujZ97FNnXqWS42o0pUkkaMxdE/cm7A62VmTt+6/4QTdCFdnpGJjX9aYjDWCwCzX
MicxGw9iW4P14uDqwI96+kYViyLQdGqTT2CCxnUdYnqMtVb2oE8xCQalAiO6zGNNsXABgQbqzlFs
29U7t4jJjUX6tfE7eNAuSgxZXvtgVZMzuoo+sclU7/PlCpLMsI8+pnf7DNXOvFm1TyVA21zFxmMf
S+SwU9Qu7rA94Ws/GoUuTF2c/Uluv4OKM5hIVVwAJCemAzcfXKKRW1ctkvQvRAS2mtqUsaG7SjxR
aIL4obdes2G/ei0EMsnhT5oGYseo223z2Al5CNeEPPaagIXhHQcWRtj37BD3V9sauoLVJ9TZ/TNe
InrrW24JClWtUgS0u9UXhcrd+8g3l94wv1cC+yOSNOp0eNTcLrBA64nfuXXp/6GxrvbCKibBk4Td
BD13Awt/mAr6GL2PONli/9/0ilNCoDzFWGaO4wZbkJC9SK/DO8OTkfrspcUbtbsWRHo5FOu7Tw1o
tbVdTVL7+8dlpEL7hTLTvrpJ2dyhINF7Ns5RwEuWkZV8XRoZaDwd3Wu5Ccyv26Nd3lZt4TXI+kj3
zuioPSV4tOxy1igKLxO4FA77VtLOgf9PUkSwuzzlbGqh4qTb8ULu67oqEA+p+6eX6Vs0N+IY6rZa
gb4UcWK3LXpTif+im6c7o/VuHYhoIvlSlFus4cwCD3J0hoePXszEHfeZjgzwNfSU62xlScoCUeqj
wsbzdITSVg02FZ4w4KIrsWQM3taW4sbPnQwGJa++wD44EAh5AI9OmYhX5ngRpXjELev8QV5WtIO0
Fcq5T8JS99CntIPfURqb0ZQCH+o7x2qpHW/+BB7+KQ1UI/z1E1hCV25T9iog9OPX1GjfoO53t+7K
T2iB6K10VKuDB93g2j0JbfSxjE5j19lJgS1SQelpZjymYaVwW029aUAIMReFfTIqrQ9fZdhbw/rE
agXZJqwDTzwB12hx9rFwNN/SKMN6I2qyOPFuzKpoyMxArQfNue0NrkuqLv/iU9ps0Yzws+sKMsgk
bdUIFsYsRLdZfT7cJzJ242vXKjx8hZTG/06NGVQ3KmjM7DztMnXqSt1QLzNajHvnK9RMu4ITdAg0
bbS3754WBFKfn/U9Qn8QcCSimm1TLYVtdNDxoVJ97D9LEqfQKglG0pQlgYZrKYPMOp18C+Tfd0/1
Lckd1cWkuGgy2DqRo2M4nL7kxbcJzbJXWjM4YzCJx0VE/Oz1aCbqPqQpigKPyEDjhlUF8ZxruQJi
VX+hmBeiPEQTJQOsFRceE5eR25cbkp0sI9an65Z2DwoF6314jf1hvu5LXOxfZP2rzmK4LKDFxHYn
mY0nMua+8LoStyYblyHMS2IcAauqpVytHa+X0FU2Y6lXU1Ja+TNKHJsoqfJ28uNsE8lCLFjHPKZ0
xiBnTGAIlq2JpWAtvduParvSaGfnpunrm1z9AqiFFRRCIPJYoegyZ1bz+pl8YgjSOct3pO0ag6uE
Af5pUrM5ZIQNcoOquDlpk39clWbuz0KSABWP3W6YHflJB1mvmn13nX1T38uLK1jNhFRUjnp+suIa
iV/EsD1R4EEfW5JcQwX6FSpfCrjYO3VZupJLn/rFYoDuzJNxRwnMPIxlp9pwMePInGaunLkH24Fi
2Ae9cj6hxFybrv823fBPZsPyYJPnYclILsAa5VAy4jWBrB1acJrYX5PvI8JErFViGl3k+mSvAtcM
1t0qx3IJQCu8xf59n82D8cHvCmmtQ5k+4wT0K2mI56B0Pc4NVJ3/qNtQBhuE36rAL7JY2Qn99CZ6
FbRBHuwX95vWJeF8mJCL30CY0nzfqHpNaTBpMjLsYBlE7W+02Hr7CMTJ8u3yddjUrpDDPJ1QHgUS
nE6gbalFsM0gv4RAJVw3ayujRgZ7bG0uOlYPlBFrQU6mXkgKRhm8uuG20jhLkKlt03C+gF0n1Ui5
moKWTz097WdpMlDi4xs8QSNc75zd2B0gFkNkcHAhrAesSjW0/GaqNLH3HZg+R8wwG6e7B80djSJ3
xd2V4XXzE6+rU0g3hicS0bGosx27bbLfnfDkt4kLpqYBv4tF0szd5k/+HusXE+bvLPxPdlR4IEJQ
H3zBfjNIA5ubfRt2z67gZxzt/62eu9G1xsFZFqKFXtv6YDYDAJ5rsQRwjTQtrDhcyKWZ+EDsMFBO
qo4CfER5D/LKHvQCmNbbv5wd5BcqhLESu9ZepmhNsA1N2W0GQ6XjWzRcRDFxjTC8TfnsAdP4tI3r
ZFhX1uIG6yUjK5V21Q81gNPtbSWxF/jhvCdmrbXJpAKYrEO9exn64yqj7yxbeQw5QCZiaNEbzdGm
umdmVmJ4rIY7d0GbFpdaQx6h6K/+qJKd8K2kX/u1dfeTqwmK33PyID4p1W9S9H2qgO+YVaKXC5Ht
Fll2qUpGD5NNSbYlFuSAqSVVSMB4J5CBKYE1fqptMHxEwxfKrXLprWaui4L4c9NlgOAhS53l+XGd
UwgaaqU6y0Ofxtz1GIBWwSUm3oH1oC74KBFBH4M7pn1EfeXZQTvLm1NH+5aPX3Ee+SplI1neYCme
QM0lBDNIzyelqakAfCeCx0Ir0bjQ11qXOe5H28oNtIEss6TXrs/+nzj70wzVQarC6traIRlO0iOv
fnd+0Xuy3+VF58hIDQgXoiTQ4IaOatizW+i3pJVV2gmmHmVXPajKGy8wkR15ulpPVMTHA2x1zpnR
sX3O0iotFdiPB3BQY+Akig1TDeD+pEft1TWDriz4SbKZyW77XN1Lj7fd+vSdEMb1oJyr4+YDju5M
FCyK7nUXTDb9QaZ85Yxi/f9+ZfwwuJbJtoBuqeNRSJHtAdWDSXC+PImE9GWGebibmOOHNd/c0sco
0q4GR3HL6iwuVwwbyfxgDubEYgRkET/qpX2/tSQ+fH2M3K7IUknAFnnrjxlxhZ4ouK7lJkqTLfmL
lYd9OYVRa212pbzT/MmzSwLTGTda8bU9u6oF8RSVZZ8CSB4jyJ1suvynnhMQv9/5JL8/onQHEu20
inWSvVd1wEQ8Q/aPiRZSFObz74ZaROKUdG1X+z7f5ETr8n7T0DNXXKRLiEDA03JvhK0GegAJYsW6
MXML4speOtICrN3EkL3HMiCohv+1/C8GAT96IMG8a0Q2MIfRgV8saxJOiRJWmBLVFTWAKz3zTELZ
R5DZCSzmiBNJZNp4nb22xl3tahOCyKb9KnLyE7vZQr3MUNbsWRifbsn1mawpNj/dQzpOBIoqFpRJ
oZMlAHGW20Ao7L2hB/9KeoAGKpijXPHxeTP38A5VtYssPTUCxiXPItSOYYdGo5AOTh6oBLcuAD20
mx93hMGJWVTeBSwyFdGX6icTbFcqwnf4qtAwpTUIE1JyEQxpz7pV/ECA3vzx38e9erE8dS6NFEHv
OHE0uo/0aSSR/x00mBDJRQCynFkypTXVqqZuBZlMZ9OhyEF3u0FnbXCyjHuBIknbzaxNgCUUcpYk
DVtMXqWDSr1rALrXiXdI2ORXnj3BJhafvIb6LOLwFzrDc88sd/OIVSezUarCF/oBhPEpsDnGQyNp
A7BAnOGXp7IgAQ/lf9JvmnSCle5yASdKtK5tNzZYz37ApWNPpWYrj8AP3aGG06auZZFG+7B3Lm+T
AlVNUPEvi5wjhmBw01a+qL3wgcW6kQ6cbhnFZZL9GyfgwZ4VS0GoDRRXDhf6yo4jKRz+eIWYGJX8
tZom0RBGFk9wiEJhcbRG8bPtwwaEmDRw30bplQFHgBQtXTf4xaEPb8ULnf7+/vZSatDYv72LzDDg
fpmAvstRO3Yi95yLKl6ZGDNEVWnqa8dPjoUPZzlS0Yg5LHG0pKoEm+zO+y6lVReGqbNPfmVeeixU
Ch4XtjaP3+k49LOUei2Aglhsm6dpiugpBvsWaaUpXDkm20aFkP4eNaIATgyrg3tPGf1Wot4RuZSr
gQtBvOcppZp5Ms4rzpM6B9rmGK4pAgww29ZCkS28yB2k0Xux6XON6DsA2mbUbbpPAJls8xD0I0t9
CQnlXunHRPPlHWN66VrmKksKiZJiIy8jRcPt6We7WrSmmT/0MMW8f4G4C+x+U6k/HTiQvlODcKz1
3Ll6G53V9vP30/xVt86ZutDO2GJv7q8OIUWNeHD1bvmbpdSFlCReIbtQE+kdE9qxhxlzl4SSLFRF
yu+STaGDD9WBCXJn26F5AO5uemiZmYaWbqDRsQZ8LSUQbUH10nec0QuP8iMrqCIxeXz/LM17SVsP
TzzAnoVgaFkinWEnTz10W/Lx/PLU0ZxEm2VCBOMKd2AMvHSEX47fWcT/gq6y+I8tgMx9Y1glKMh/
0+q0MGKcSjDZKZvSRcyt8KLz+uAAsvAeHh8Hu4VEYv+2yLiLLK0NcOs9InuexVZuF5MgMhB1pwEh
ADkV/SvB1JCA301+5cVBTyIafoYhwBRF/pR2NcExjeJxvNLC4vPZ0lpe8wwDuuyV04PP5O6tO0ct
CgpkYcL1HEmlmmthQZeASVtIQuobXjt5akL4hBabtZ/egQH46aru6HLncpKy/dXBgau6X4d2A04K
aGDPJTGgjFKdOyev2Qbf1tCVPn6caQ9xBJeruZzW8XHA92lLsS6xJuXmnJSCUJAnGDf6CtTAkzYZ
RVOf7kV5cE9E2Lh/bqSBsyJqLeIZbM/nvYL63y4IPjO1CzRt29zdj0WHSXiXHCo7el2oThTdqEkE
S4+uYQxptu74uyoiDboJ45OcR5rdHjZIcFDfa2H0RpqX4JHYHo/SHNg2O3GKSGLErGuN5ANkIGgr
B4rRwq3wvB6rMrwqwxLayM/YddRVyePECgPhRTR+KlmMIBJnlCorP4XzWureHy9Vg9bGPgfuCOVM
7zKhBMq8nz911UAhImeUbOkkXkvzdhwqYj56iJjV1hBfPoVD+zQYAFgHaiQY+PKdt+KeuhF+qpxi
A9E48zMzxgfOvFM+qm6lMNqjgdcm8u9piM3F+ofNDq8GFQo6+tlL3ydzbXzWX/Ur/2x0uG0dJs6a
1yU13i+Dh21S+lJTxueoW2f11t98jX3zEHZdtL1PDa+rAqs7dcQi/wPV9obr0oAzrZ8x43CopXZu
ZeLWn2rfQDuyXP9Zwzk8j9P+8ypp/X3ykb0FGmhmJ3CmRUfgyHEr7wRYUbWrB7xWUVqFcY9Z0TmB
gxVlQF2YxAwCdnQK6rerdHzMRhWLpGg3qLQsVGr03BQMslsR6PyUXirGVDZcLw1NCnVcO8JDvuwm
4iL27Bl+4Cs/6KEYTCstBU6mUc3nRE8cWKlsYb3EhxfMCMtk4ZmFn02wU1bZMfEMjIT4fWGtk54q
3TWYwUZ0TJMaTasVx/n16oWhf93oSARniND5XjUB/Cqb1DYljhPftcwfQ+yBv11S5vsggwlPZjdR
9AIBNUcfxzkojAaaKkxtLg6ufi7m/a1tYrikJjLJ+ItiucO2joXzitdW2QeBwAufwT7c3+Yd0rSC
g00DABmZzHOsDkJQxz8nYzKGxGRW8f3HIBW6CcWa2gkx6w4/DXuxzisqjv361RGUJsRqW9zQMbnf
qznIGpNqtFGweqg+Wh7mFDGLYjsBi+jS+XxW4eN9PDiyy3TZk/T/bY2IxCbUEdQ5Crd8OD4oQR/q
2MHTMXyxzQDDusjTAD5RjVopRJbq7mEntHLKOOWeKK7YMjGjhiMcj5d9O1rJhIHdOE3aDTXzZeBV
ttQuqQ2TNxy7srFyaWznNlrzuLVmDwbi6iSRA5ADs/GracdFZl8ezzMnIGwRQ029T+H4FEe2N5Uk
kt3tof+/y8XLAzfeG9xYgN2I/yANVhRJ6atdxHuSkfzj4aahyeVJopVGA2V5IGG+m58/QsZvbDBP
3SKIHGIO8AxKnJmNuOFRaK7QU2Pmoi4buKSR+w3YOTRGY0SlgSh5GJGEs8bcwN+4QRC9Yysg5SC5
c5wV5X2hpMrpkv+SUXIKkPs6O1Ajqz5+wzbJW4FeYGacXl1OsO3PgjfCUnralSMJu+KwckQCVjdT
0WSK1nhvySMKOm8KWwwa6/W/mfVB94bmAq/aYRMg4MSqcyiHpldgo8C0HDH0jQ8opYHffwnQx9IG
ZaF9R+0bXfE9w6Hh6DHplhJocdUj31lOT5veEDFbtRoGhJQMjOMcMIh6SYbq6AfAGnJq8CShJ9QO
jtPVC4TnPzJLYuGmuu1FtqaU7TOHVoQQQpRLt9/JqzifKrGJ2P4IDLZCJJolQiSiLCh7AmKtPhk7
gl1wfU/xi5UIrJKpX1Z8ySPoToinIc2EFh0/Ueedbi9maig/du7TMPYp/sFBoj1HHbr9AX0uWsqA
SNTY9EgmJQNT2qJoDoDOi8XD12Rp4MInJu/DurCaenTo65ZrHgngCaNpd8Ji4NuDZ1Rvdx0TXF7C
/5GY3OYG+uUaNnXC8/4LkgcY3/CPF0v91OLxImsSt8BP8W54aWEZkiKbryd31BgcdVL8hD/VFrGA
11Xo20gx5eo2qRaCED0KOLSd4mB2fei/BXdDJUmZbJktUt0NsuiHrT2+Mvqq7BrH/sts6SyDmtNG
cFrVEBCKDqjzoHPvUmHOoGWxCZhPYJ4s8Iqxxe7LsfO7EMudsnuCOdvNocPaffKOBdfMASZKjss+
kOIQcQzB/Qnnq7R2L3TssZZyb2BOvH/P2SnY1r23GK+hGdFE+uI79IADbhKac63FbMsVJqCt6tV9
vC/wZDxl4tKEbhBXANASVOSDdcLSAuEmbzOQMG7pVCIziL29WiXvHYU+xoq/5yCKwNo3uTi53+aW
2PJuLtYLMoOQPHFcABlmvGMHypDOXuhak01loGKAMTWLD+kmJAG9XYgeI8NH0Ah/OnHgDyT7N+IA
xTiIJlDrm3hm+SK5a3iYfCDImxBinIje4V9WAdTVVdHYjnAlRBAfUpOzCbhimfqlkbg5IHALLRFL
/YGoxVZmTs6Inf7YXFix3p5gfid7QAGPRCbMhNIpAMDSXOPwyR2+Y+nX2VcWmyZDwaH/LKR81ksJ
CqgqYXHaIfAUaqmLuOuE+gkQEBDXfP16/g1LBuOgNkC8T/d9K8DpVrx7otrvdjD2w7YOuUyICXW3
TX3Kw1brh5YA48KaoFFVSb8XC9/xHSN/v0O7uWTI3sNLP8OMRb1tl9nq1QpCvBo47cXOqaXcJhxI
GbAS4yJLSNX2GOiCxjjQ+5iLzD+nfZsI86GvYsqcdyJSPF+ieq+SmfnnBqyGe5OdNG/M9HQD+12m
AFmg75hnyXInKtZiDmRwuRD+K1e5WPd7Sl/HrkNSXf6LhbwKzvMxTqI/12QgVqe5dg7pk6yqrQVb
/Ncrm0R+ASZdXVQTN2FR9qS0TumYO6K656xwEx38sHwC4NrKm+q/EmkehuzfE5IGNsDysmKBXtj9
nlfR8oxHBMZZqb1nDRUVCJFmawqyXxVn1+RuQgvXK2UhcSAPWDOjmpKl28LriMC+ryBKYGYqCAFi
fhqBYhLedlkBgSkuDBizOeg9wFvrVjtzXz58XW+7IHh+v3Xcgpseuxf87Q9foqgoiytDBy6X00RR
C7SKZlvWbv+JM2EeUuF7bWQqjhC3qxN4oQbLU59ELb9Ld63DTUS1ajKF8p9LUWzNMBey/1YTms0Z
yckOwY3hn0k9Zwiap7O5YgqS2yow85CTv5+6vFtgKsSZvsn4zN6mgd0JUUSdCXeP5zOTn+M7vC79
t2mf15DLbLhXlDHmqEAUTAA0TP7+A9OvBL66nlobFe/iuPc7Si3T6p8hMTxKyaiWPt8mlc51CB8I
ew9RHxsc5wbHySCZK1KMjMJz/0XQm2scPpvSh09gsqsOP4FDlnADA226HSHSJRXgs93nAKP7BHTR
PtLjPRZf8IwTY+rM4aeuGlz9dZMOQsAXB60oCoRQl20+lwMi2TS1SVv/eIQMV3u4o0JsJvbv4STx
DaQ9/EkuDVy3PAEFeJhqaDxBC/0Rtnqj4r/6qZi5IK9eVPsCmn30kHebFVvYTq9Gmss5GOta4Qfr
imMpzlRPkgOL0MTwEaFXm4OOVowtlLfBYNjjOnbc2uOGa6mkwiHB0xgHuaYk1sTQGHfUlswnMlQz
eNXx4BHbgqo/q1f6eplgoY9Z/5Kq/r9bkDbZAKcWEAFJQvvfaJpS7Jcf37EDBKcPo6k9wuxZXydF
i2ZPFRxp7UdJOkPvjOHLS1qJKoBsRb3fTNsU5ZHBjIPn1F48P6KUZ7dyI/HWw1FTKxrP3JZ4XROt
GnAv0oCFFSMdoZ4fPMAU0V32gQaVNyp15LsUfzcYqLcSWeOgrdU2OqOG0MSuwUdeJp33XWW8YZuj
iP52A4avEXJJOSK/qqTUFShqpxMBetPZwPLaWIh/sUyW0sNyQRkTdKAE5sGFltACybu/FsI7/ZN1
o/7XeXlAFEon2kT2kuMSxz9/31/Fklhd7YDtEUZGWohSS1L/EJHHold55oA5312F5hwcr8QYYS6l
++vDti0OQA8UqdqeMzlrsJXZbPGR8nyW5ZF9zMvuUQjbmm5RE4IA6QP1JyTeGd4SJYMVNpvh9zHm
euD+ShKQ4gqRuoerrsh6oae4DubwATqKTlhhIoWtmKyVQC1l7Do/1VGvBWbvK5RcxE8rJaC/0IiB
7CgZrniFjAyV/sXDOAiTDk28zww/9i/ouB6FMtPksEiEmXR6B7qbgwnd8b7oPwIP0u1a577p4FWU
Z19erue4tQ1GJyY2nf89L4RuejAtLmBlvjAf1xP7ohF0I22n1IyK++/AUm0D2eS2UXahnwUpplv6
rPWHzhLuBo5CZu+2/0Klw4Eb0553fgCsJarQQkqks00fBREbK0tV1g/VWqfB8lYZmb6GUUEQ3OWo
+lSwbCb+Wt++d7gY2OLGT4/NTfPRn6U0ptfnkV7n3fOdBo/3A2Ie38nZOJpgvOCy8h7XSNJiyJNx
KGOT9yaoFw64cCjVfQSEYXrb4+3uOHtKir9M6htILfMCaJy8G86QEYOSGKhC4KPOQFpW1D9NZLfD
AMa2fh24pkl5MOnE7w08BTKA5cjByiS1yrQ0PhymucT93uqPCgsSjMGK1xTCQFFNfgod3xipZyNy
xUu4r6qMMSSCXlJjZdK5/+qRN8s31SPDlG5BBi3gqx/OuTOA7poB6eTOzQDHud63QiCiySlWc1/8
E+ppcdm8nQleRWoF4rcfN6eXWtEnzT24/L9DldZWUa7iQMwyVED5Hx9dFuM2Yq6RK+JFYqLoOOCY
wlp3VA7F1nM3Nn8i3LMZA35UnnJLSW0U5inT2u0TKMD7upJW5nS+8DhrbLgHCBJKIrW0AiQRQKSy
O7By7sTHVez0f2bCEXiO4E63llHdu9V8if+2dNXvDklrfaPrIAV1o9rI56q7z3FYAxIjthMneacQ
Pj/qhOiRn4DAgYidrQbglePxmTZy3WL2va33Egw3QTj9QlTf08u+iX28VuUnzciXlC8RPUPkeIpV
hMUkGgNxqdsJZwfVaPDxP5SGkWhOZJVzcJeaXvN1K55U7VipM7il3vJn2/wihVAOJouDK1yZDzpa
47zC7GBOHeSUp1OYsaLsvly3ZV7WdurpPm2CZq9+k+pjych0o/6swHZkmOk7/HoYufL5dXD2lqQG
QCFqwxb9/06JOWQDS6uCFbK+JHrpz4D1I9uEaPNgq0wMVTLR3LLXUah0HHJA5/pQ20heSfoFJg4H
FYdDuKndNsk2Rfut0uPheT7/l0u14IQM3oQS7NgAA4VvnOqvngCdyP2TwCPCtbpPWjBO/7XyecFJ
NZsyukPuyndjsZuIQNysPE2HFoPVs1vXNqN7ku6zpJhalbxS08oLD4nRM8jgG21Z4NO8K+H+SeP8
CIIasXfLFAxTIwcGLE9cndvO9Dkob2XC7P4dMANMqe/1MQENgBY3qkBsezHT2SNyJ9k3Ax427jLD
OYXAbq8oke6OHU7AFXlGlMDClJbBts2dfcp2YCxbvYB6b2jaLl4NJK/J9jnm5ytJjlYCxQjVLbQL
gxlNIyGrnMuOw9uNMuYRnhGr/SKk9KHu54LtizBhkrwWOEJFqyUOpu7QW96ScvTLfhwSI8pVoIW2
ZND38tvZnAEesPOmfHHYq0gGYVACGGk6GJ2Owkwg8CUnRrKSEM8H1MoOw7cQZqSO88IKHMN32rS4
2kfzQ/HxuWM+R8Wx11JVhq7KZVoCUTyEwiFrKMn7jU1/k0iR87peOSF3W/jOgOQSLteAT19Eni6l
6LJLao20JdW9Hz8XtSgXvZM+uE+HJFhr3FYOBg6MHbrbVY7JXLPCeGADn+RZPUMwzu8EemX14116
wbCCb95odpBA0YrVNHAq/3kwxRA/SABZ3vxNeHtkyNrUEqKpfLAYTJxLGlhqIlRiyPVD18yomapi
13QDoiYQVhEekkNCjBXfgGJtk8caNRwYpVPWzXof5W+6FdTukOF+H+3ArR0z3Ljp+SUjEeQVFNeA
I/zVnCpkrBJnJTA2vCwJiXIF2k/JnXPQccGGY5VrgS8a/fg1nz7FvRv52eBxNjJc0pvvUxEDNjLt
Ai8m01aTFaapg/QN1uxtapf5WpCyZ5gCHhMOgrN4LPS9VhZ27TGwkjv98d+r+qvOlWRef7Ed/VMG
WfX+Ihwai+smDYE9pxe8a039arA5eGFk8yEvCLZONN3QLGlj3lQIHPLGcPQ0UPmXwZATcgUYPazh
Jq8Sj5+5iPSOVMYZ4M+ksr9JOw/lWzGG6Z5TtoO7TnJTdiyy/zPN5qQSn6mNk8R0Qr17VP8YQD2c
TxrxItn26w8/9ra9jVMyK8SnKgsZCODdGUEdZY5j93aErAIqGXx0vqxacdNYes9/mptZv6hm/Ly8
nOq7WKiWVHzh1Ld2JUM/JFyA+twxpvwMQ+8mKj6I5omSc47SfwvutW/Mxf/97zFaq0Gy7q/jDqcZ
F5Stchc4Mv0gQZXR8iWbc5gyBTVd/rdehuunE+vLGZQ6278KbFI5D+p6F/HF3S+SNdJieKcHTj82
r/TxEZdxC9ZMzI2E/QkS3rgDAdTzndqc49KqHMpx+FH7q7QVpt6HyR2cCseoXduJcIjVryrEjSvg
/YOlzsTWc7xjZQPrVAvst2PPvPTE1QvlZ54U7tPixWJf/JZen/1YfV1uAbalrziC0lR013prtU2N
Oq89nV9xdgp0OvCKReDgoyOMB5Km7X48rSrz69d3Ke0rEyvrotJKy/ARhwtOg6642ecbMFG/hNpt
6wsjld4GYaW3JJ/JKSvMdiIol6P4xovxV4qkuzJERimS7fQaxhFVM/nsTm+PpboL9LZcAf9Vg4y5
LHq7ZfrdilzkXW8yYG4bSQRB4qWEWQt34rCUgqLMIQyaESIWOJJzAe82iJ7ZpASX8lLdHbLF/FdG
nzf4E6tdP3C0h75VUjx/PryyQookjvLBlzsyC7ise/l74ijwAdyFZ/eMZgPX0hXCboaKFSE9wtxq
JDv6N0pFKv8dUDhTlTaYug1LWYN8Ctsi+c4HgNLsKnjVAEb55sFqHVWikFgC64N/bM37DCVcAfge
PzKpFRO63mIHVs65kCclAd0D4cIq6hDuKbT5qvuZGcZ/1o0TP11IclK64amBcIMuy1GHHoXrVVUM
WwBlDuAWGkiHitdj9NFtAXfhf/emrrpHbIVioLm24zN3OH5LQPNjU40uR+ERBkF8Erh01ATATaYz
q6i85SgNeO5nFT9NzHSpOSHjyVQiCc9TdylYC1WAEuhdDZFmDlpEwJDDRZpJBBwHMqGcUN71uRml
PY4h+2cQEntRp1ObXTeppmP3EgatxjrywZGM53ioJv0liqcNrMCDPAugnFdcv35n8inGYrpG+3DL
M+dFOCA52NxhXjL7Z9jqtAEgCvphMiKilChA1SoAeM+ZQ6qIXkuL3jIDgeTQQM2OYoz2yyAV63TU
kHvQVHUenUu0+9J0MRL5o60EldbAAFx1oM/fZbWR/+zIEdFBWYlqqgUbGYqBLTfN4dzz9FIuBmFk
Ezw/tzDIbqThci1rn0dhABqGhIqhQVTz9TB9tABLDySM8t6I+yfyGIHWpbpf9w/XP2OYdXQtyCt6
esd1455dp3oeBrtPB7yrFRStJNkRrzxRj2vtOhtjJnsfPe8E/8y0vlIiEFz/z73q91vQhimQmODC
d1pWkaT35K6DVjQ6i7Pbtna2wWvFT3ctTeybrdYjMWEzQBt3+FpR1sidfEo+w/F2yNHcGj5FdOd4
v4+cLfHJTBRObUInnhlwIGVuaRx4DklLcL3ufJpip/GweVeAJ/VIhD8jxBGq+f6iHO4MTMNitnDe
wNNwlnmXBi4IWZCA7sRs+TX6ULko4m2n3ctnpZitbF/vtxIDcPo6Nd/qdY2edU6JvoHJ/wz283KM
ZSVDUM4v7vpa1eBgjMOSQ/rDOHkTAJOJcrhJecRqdmm0l3IjWNhtGkj/frl6LEwoFzTsjA6HH3LF
PsDRPPg/f+wT8Heum6MC6xyCVO1yCiwdswiqc2cr91UB2YBp9TV06GCr/pG94pFbSYhDrC6zrQlM
4+Oz3n0pRoUc8DC+Ep2HfBBi8OXVSujxwtHApiqLjpdUBkXnETmOv38BVOy2qJo/GBullwe+JvJ4
VxyDPXTm0nkK6UwYM+m+spmzIbexpfXZk/0/6G1YDkCSGqc0vaIXTuounIV2/79cUrb76vvtqZzd
8UniENXSsoFX1AldyxqnnQ64sMaVsAWJHZeRq+3jN/i8nAE/pchM8SPnQyqEwiaOGl3vcFg5frVe
GAZQUyvFP/gWC2Ubvxa9Je56Q2NGlF2QuyxlgxI8VuilVuoiFQD2X1/LUBCTwCq6OjlhTVRts6LP
pRI2C4ZgZDKc3fH7/gx0lkoQOXVUUfOpnRoU3+4uWIWcI4gRP3S1lxrXv680JXX69KicQHIuJj4a
a40m2jtGEdhF+amrDVaG+4sFh2Dl3PbMs8jbFbBc14PKm77FwSsyOnwD6Dl4qJs1k+oHsW3lI81W
+15yQC7gnbdSSXxLmwtx1cgqCFdW2AfUzo7k/aepL2JWHc9SuOqQ97FV8GdmgbQL1XNzI2g7rE7C
JouS10JkHvOwDwaI2xNRT5B60XQs9eECJWSanxTbUFGN4yBaYORfGCUxRq72Bq3Cy/C7Nzor7alG
vSl23Yrmst6YSXMgpt0PRer9V8HM01SPTWL32n1EFTFo2jKjnU+FN72cqKQ8YEspqrFL1heJ+llA
e1aFUZTIHhwticeKGuDOL11lFp7mSg+8LXVM3cXBWGrwfk0aWOo2Q63QmezKJpdqn+q/f0usxte8
AF2Ey7If3UYoU/BgqVDnwsx1g3BE1UoEO4BFGnZ8WRa/PjJUp5k5JMOw4PWPVOEzIW4XkqP5st3F
ho2JI1BvZyu7ov3QYuqSTzpNKemnxals0RNZRo8euDzcryptWjJ3r6NdshUdJ78/pV47zNWCyOks
zA++zoD7EXpDQ0IXLoD/ed68vxsha8CWdKH4dGDo//XCW3aFd5fx8a99fsw+UuLYynj6eUUVJ37q
8LFLFK/EFtH5lnZ6U4Oi9Bb4slO5nmbtOAPjFgaDpjuINCEVsXz9NwhqDLCDCjll7PPL1rJGM3kR
1FxzbFK1tiIQekWHd6bMPzDiYRNLblanxB74tVIxX8NrfyG/2FAUduYgX5d8vED+liyHSecGJ4xz
YVMnkI4xd1iRLTUOH/3hRCvN+S9XiPDZ6ZgUa8pmCrXjTiq0tBEAdOzNbV9PYCkByKFw1lFkCmgy
RYgcYFhSPj9WLKHrEeX9OT0FE4/D5XFE7aGyFD3O/3z9K5/SmZcE1oOat2O25hYm8MOCht184TTP
QVg0gC6t/rbfs8NFdD/MAUp+oyfYz3qPkMMMW8uodNGtGED5Nalrj59exI75qFC8PmDCsQaJwbw0
Z/JX2+SMMHlhbU+1MQ7YGpnNh8v/7bKXn65oVODbGZBBJ5qUrASQuIXBAlXVGpkwoLA2MYpn7GYx
Mj+WCeaO2oL6km8hWNHMWwOEKyz9/OedHOEmO4J7OUnBKbVhXiGSkLTFr9y82pylgjqpXaykYYeu
/FfQoeQaGsFL4Nhik8rJ+jCvYJMAMNzoOA6JfisqREVSnhYQOaM0Su8GazIJP04WSfLYuIU0cxdu
tdjEOOLGvqguCMu8O/d37QVIbrMGS+yt7hqM5aOiCQw6djI1e1n0jiBVqEF+NFKmZ3iUxzgz7L0y
De/VYZJHwJGxUvKSJSjbcEL9NIXA/KISCSlHNpt1GklM4SntioBOZTwz/TeqHNyw6xSX6gMF+hnD
epOQAjTs7xuM0Ml/MHeAjECm7RFX8PZNOnyGbRXVJ6xAQrbnA+NZozgfkPJeQd3LOG/tU7ErUQJv
7IZ62fN3MtQa72esI49al76Dc4lKWtHNwEXxuRIf5jskRFNWAA8v+ns28pI5rTKGp8vH9luEWTgJ
vE4xSj0CNNXy/6jA/iD4TqVIKD+dD9XFGpgmg4qn0cbisBdZdHkJ739iJvEqGudFRh5n6cdiSwP8
djkr+SNXAFrXj5rMdwi8221Bz+IUb910xpYEmhdCPOGFpMgnE8NF6tuO1OpTp5S+EDqGbydixs9Q
9jzkgNQeRONiD3K9jU/ENdXtTtESciOFwGgl7cQmBV0PnHyAZVRy9+eTVxfzqlCMPsWZ0UdE+GbW
aOu0eNG2Y0hbPHXksDeqS2JkzyQDxm2LL1ftMsDRzq9EeXMppevOeSAFB24UtYFR0j5lViGnhm8d
VKzrQpPRs+v1FszMMrrVayMOElTmWcgEBaPGKyRlcA7qviuzF0davs8mr8bC3cZB6pV6YMnA+9b4
EMRdX8ljj3iE8xFW8Wl1GBhg/tdeNGnWdI3VxhdHVIcw7kWKC98Um5WIbUtm5dtQ172yi/ULm6zR
eH2ImNB/AXE7L7ZnDiI2HpmtyhzABpSPvJIvtPcZSFgRshjobjNBZ4zihZGkTvYZTotlesCEMOse
2zSagvO+DFd0MAXgA3mcAzM/w0n9BZoXLxHVPeQGOkJERZMpJQ9goIgVFNoPIkWX7fj6sr1FAPTQ
0ovfKWCeiYl7w7AoE+N7104larUkf8X2vJ4v4jdzM9mBVaAUQKu56LsYbMVHN4CQ/B1iV3R4Uu/D
DTVFxpML/K6sxdG1EhGm3uVcDd+e/AItpFjXdqeJPC0TI91Kgb0U47yG1agIXXvkxwqLyNnE9kIV
DEL37kI3DCphRHIguM9okMQWjrkBLD3fie1UyPhj5cCrjnHYWSrnzu+NRT+R59vDPKexkF/Mk2Al
H1X+Ls8BMdiPPbnVZHh+MWJs7P92dh1YZ0+a9mOcqNNxLEnDqNABypmxNwsqaqiLpFj5+DmANGGk
OgpqLfU3B3snVQGh3K8sQdUxyMN4T8qPmkBzAzO0c5W2qWRyp8arTPTsGoXyzT81lCIbnyDIraMS
FTz3uJICQ37VWrpGy0ZVEbih0xRSiXKTlLMqTZzlUYTqT55aSungTDbEHP6OzFkc7GvfSIP1LS2J
y41LER1gXgArfOhVVeb15/MFQTCgyEYRR+6TDT9nojLn4jaVApvkpm2kWTPVMiml98Ovz8ZBOHgI
BzYflZzBvCuz1MF2Bj0/2yDSTKHF5gJmtnfsMLqoKWHd39Xg5txiRMw7t02u7wYWcQ+87HTnL6d6
t8oS1OOZG9nlsiAGINw3vE4rBTiWEWrBmetG4PD/OXt7Tk92O1do/jcULvNDMhZX3lNSttdpG+qS
4cqFRK/7SB/YF7Z7eizCBxXNvNrwWoT4wHUBVXaO4bI+v21yCi3EhLC9GSMATH4HJ9TTfvWZ+cgP
UF9qRwBEIA51isfelyoT+uLhRMOmL45+1f0aPxOALa5HiAfdkq6U1sB+JKGHDcfZK9KIhe2abE4i
0ACjOTZzRGDsxtdGgOglpqVrqeW/nHkerVplEMO+Qmu/iEhF4hpFzks2G0D+iNhDw34Qw6U/giox
GzbXXT3vLlAPec3grAibVNhsteiDQvxUvMRsGODIk59TYItw26mSlb1BMPmoesj2YmnpQ8To4F2w
D7S030VP8jiSrQooutwRrTVP67AUkuwuAztCqBRpNZCjYHHm8dsvhaZTToPjJPAp7VyydAy+3Pm5
cZI6afFaM5eSVBiUc594yAcyBTSJStOZ2cdRY0ZFm8IWP1+Y7aHElpenBf/MD5KDmXRt7p5F01MT
RoIQuINR6n3WW3jg4M1ZoVe8XHUzZeCSytNw+7B5nB3HV9gKSc1ajj70V4rYZAK6vDrarjD9cYnd
M1nYLDWoAG8bneWkwqKQrKf57cA3FU3AK+kPZdp+OtKEHX7CTRjy2rPA/YZYdDPL4frWvN/Qjp4s
Zmp7r02NoqV8AZ6Rj9cms+heyTeHmXUe6boJCUlThwEv61ePQdWO+OrnYaxH4dkgGDDZZa4G1Z/M
KZfhsg/pNIhZmhVwrsimVSK1GgTlNf/lOHE3XaHdVMQ9F4Z1Sjs+mfDyRsP1OQKNbqBRm+lL53BB
6+nz2EztsQAyJ7jgyACjfVADrK+9zBIn7ABrIW6M03ZOZjd97v/mGL53fzcNSsT1LtljL8Fa5L5L
qjj/btyc8fwJzFpHyHh+k+xiuowMS02Qf0suyO8Cahz7ozrMuPCotNWuetqKFcWkCp5MrMGN74fV
q/IUq7FdxvT8drl+7TdiQ5U8xbw8t0Mp0nAEDsQYIJcjTiBhWs58GOvlR7MjQfh8JzbN0E2gVIPA
F125zDSkPAbFnY0sDfT+06WV9fJvbaDWkir0otB4ut7EYSlEJDRFauCkge2zQqOc6B7kyJHlvA30
lgh+BMNgA++03frjfECOL0SMksBXH2HyTGeCUq86D2MsAIAg6K3znej8wG+v51ShoCyiSGDsJKT/
OpjAD0SZbXS/p3BmrgHpEc6TlkgFZAG1Tp60vpTK5WB9BU6RKC10tbeiwNI2S5aLFf11279v+FqB
PXjvnKfJDdjqMFvSD0ZoFjECwFVrkK2rrFy4g8e26wzXzSerY7eg8f+aYf4mRmF/wE9mU8qsJp3v
uNqy0YLmTOqq2wD1M5Aod7m5Zpx/DHkhgPRM5TrTz+D30AT82pC6uR2OSSAuHw7KKOzPa1Rkpgfn
8yBbx89dn49hPd3xVNeHLt6MEVq5WZ9FPqBEvP4K32bo96c2p6QS5bRRPz/X6FZN1Bnd1dKZv4Cp
akS4Pz/kPhL41ij5I54ZFeaeqkmdoyp7FKkleypw9XjG1o/JGS2Z6dZbXWAY/y3JF6J8cFvdKaAt
rv3fG2gAlPf9BFHXKaPEldQF8XWP4aJQlMAl5mzVuv5GMZWFIGoZA005nviCRen3Yzu8utqALTTf
jBPKwRqzWE/vKQBZQjUMWfvTKh2SCCcf0FevPgD7sEEKzMBo3MgZQ7WwkotrUDc6IQT5A4W3E/NY
abxYJOS3dBuE24ptawg00n/5L34y+oyLLpe7ybPMAb+Gfh7X3VpAst8zucvIULtt2grXItyTfWTu
V9bcd1D8g9Ws30QhlJaMNTM1/dNBMqm83PiN6BFapV3NHvLfLDXKNeYPMOADDNBvBrDycza1fJOl
YHuYlJa5W7hi8bLuEQxYk6/W7+k49mWsPqVKCzY7VrIpsThQR6fJKHYpNyWhduydq2zSAkTxgi2Z
5vy5ve+ILA5T4FPoyRT+MQiQFNchwI0P8Fcb6SpWtl3zekrw7wT8198jmuXDcBVALY2MLsR4h94Q
eT2QV6W9Uwa1U7gmC4NT0WwGv1M3praorfZQXk9UPcUmMBzi+Hf5nGtj8emEartHydtqEndjVMSa
W3v9RJq/73oCTUKdtqInYetYSq1eU5BtVPLBHL2m3Vx6btyBKo5tV73VoPVyU1qQDLoTpZ0oyeXM
enJzl6Qiq0gTmjLIImw/9C52A/WlyyUj5TG4Z3NhyrXt5/U6cRqQd+RjTOd9PmPEu8x8BRrg9Ux2
CPoNucGZiX6TTVR2uk4PN0VqS7+TM07ARO+vltc+hOd0caFrQFoFzH4O4rurfvnbqDgxlVsF6Awo
qh6hn4SPhLFtQsG36xN+Kv/DwwMvQrYxQpWi7qPbEVfBQwSNTvwUi1CeTn3qzBdZGefnZP2zGhlx
ZsCBALr/gpDs8OnhG9MtFSNWCS40qqGQDDerfwwhx2nuSh8MyKSjKkdwo6Pgon4oLfUJCjiBzWTa
/+jliRWpp/LgF1ysHDTm+Lk2Z0mJwWw8ahQbVd8hxl1Oz/sv2Wj7Rx50GYu4ztfj+04EucL0yxqw
Mes9Ck5ncHHk+kziZ9SKdu7qr7h85TkFvW/vzrOkO+ufumWPRpQ8y2sVXp4/p0fgbzAyyKUgMgxD
lShFaNIPl3hN921kvC05WlHKLcaVYXpI0U92rQ3PyylV9lYfQh7nURjeWeFzFcUM/JJ8y5EE74LL
L6K4D9WnJn2AlX5ve5ZDH1SDT8QmwAHVQapH1l7mpdOOa/xCqM9+bO691C4gGVMS3j8nzzXJNE0L
tipvk2r0Xi7AvJ/Bl5K9BXA/2AB0agBRLSFNN+3QUNblcRhQ9B5FAAPvQlrkwJUq09BD1fvd8mn6
UpUxwmGkL2EpzNxkXEuPz1mfxItAQgU/cuR6Fx/rMvRQtvXAcqdP56KKPyMmhCK9XqErmzPrZSU6
An0z9sI5I+WHSXlGggNXB1QNe3Ph6TwRSsHMebb1njrEvf490GeXwlfm0N2QTgUhAKV1hjWDveEu
+lXGuJNbK0Ni+G4JOYsnsBYPDOWkn2IJ88B7lrqr2f41wpLvnNw8oicOGsH6027eSQ1rKnj4kq3P
hFiECU/wbZIunS4sZu6D8qCX0cLhNW3cwGNQ7b0qUv8udebMMj3847XYjkaNCmTeAq+LjKfhx4sq
TH8HzC9JFVO4XF9Wdz8vbvjnstWZDKhhTF85q2bluwc9WOqzF59s25f4L78L1+eqFea+Kfatp62H
1+Q65F5LmdDGUGYpSU+t5V5Jo6SM5SNLQBGJS9iRF7cMAS+URU7ffyqmxK6zVLI8j8e84BTvQ+1P
JpTWEjXbgKR3PzyJfJe+KPfND4CPmmjAh7XkaQPGYyWF6D62rFZJio3s+O7Q1fC0hwCEO+q5TnZK
o0mnX0mMOC5WJTgy7MRHla+2QNmwqTeYTnPxF1tOU6g9q2pMZhaMHr7/Zm7vtY/sq7Ob4mQ8j6xJ
TU6vyA9SkJIQcT8KxsFhem6e6aCjmuNnaLmTBfwflhSt6Oo2Vr5XUT6CS6eoZIy7/jzF0CCeVMzG
Mt2N8ktksAdC6iWZYvLFF5RcoEqAvv+Gcpg6ohuuF7auesO4BquQ1m7afCLFMJAiMUHk9085MsZx
0gAJxjLhl7mYL6UMULHHapZevymi+9s/CRBH1HYd/NsZcPLiVTjYPvQusGl+NDWIaov6HhDVhWky
DX3XYznMFOFUyd3y8AuJ0YgVgHAl7sha+xOG76A5MRB+kNjwNcD2Mk13MxenkwWCsQRwU5gSM/C6
BHpeMEsfRE3gYyvPBisKwMGgQiNr2Y6rLnfLY/hjun5W5tcbKoqpntI1Mi4GWwdMF0SSA3K1oLqD
WXTS3bvYlEIVbgqpoRp+p7CfpfKvJgOxcafp3AXsr2AhdFdphs3Vp6SX3BRR+fIk8jsAqWw/9h/w
+QJINm2X91DQKI75L7VQMBiisGQogzfwOdf5IrxZXBzpuodMjICpfqNDgPyRc5samoolPBoQXvUP
7kXEdHb61/wI2qTKKDoxDTE3Cg5wmUrpmqoFmJNQN9ZKKc0kbjpOgmnYyJ57p29LdXEN7KTRZJn3
FD9qxpyNvpNYj67eVaTypUnbShOt9boKJ/1GQ/Aj11LD3ecB7ooeB2kPYVZzB6rzVrsoym2+7oH3
1SeN7uh3jgqYGYRt5eA51qlXE4kXWOl2iBVb79Hgbah/oToQlh09+og1aSl6nngW6gytvpsdXYZv
/gMilo66mEN7Cq0X0hGAjDJXh1klVqfqLjZj95QcZEJvm0xvV4jCAWfMVAJfaOuNxuVvBrLOU4L2
UHvYPBU+kp+z2ezYWxfh5leDzj2iWdHdUUrc2A/HBPmMQVdBr7ZEtcrrqr6zrNLjjH4pPyBmhSlp
TPZkoy8L9oB45/iC2xRYbxShCJDV2Z7u+IpfXhJ6AonG/qPnkkPfumpIMaPk8AV2N2ucnyHJzU6g
wxBu6TnxSJRcU9LMnak4IuHwu8GKMycGmMYYdeUf36OeFdE3BPq9J5xNbu/LpJC3hO0GYYsKfcp6
5St5mGDbuG+T669AWmEQOLxj+gyaCvfUUr7nGehfit5rpWcjXQtKIUDo8Nl59O9fH1SuIeXulCf8
r0Yov2etV4ovkjRYtBTDW+FMWs1bt88vLU0ADtfN8NOkHNR+rue0lRcbhCt8Sj7CBdPdWgDL8IpI
Uxv4PZg2IUsGf3+1Q0zCNuFpnKhw2ZGWrFe+Qda6MYYtC+U/6jYlfUpp6kD42kW7qhDeiaKJ7n94
e9y9gWXnE+QxEXwg7qOb5WweQS4Vu1RGto+JCMhfIARWabTUp6bUNa709Si1leSXanhAYw9RQ7b+
ALB7i7bzO5usiA15CCRGRadpzKW3v60ZcIMV+GD8DalXMhBgMvc+Hn++a5ufInLSUMt1Zt/VcrUi
zo1NlkaDXUrW41nYQW86AIJcwM2vARzHbgvdqALrC2LTyO+RVQIccwWl85E69qBJuASolDkklqUa
NuDLeMx7oBXZS/JiNGpLptt1VhBdyQ9QgYREK/cZ3++GoHz8Wqy25t2XhIb8h7B4T9mhmhnbBELK
CVcdKZd608i5QY1BAEDvojRD+B73dzU+ekcapm3U33JwoHof+oSVau7hAQ1nPoi0P9rraizfRK6D
ci6TSRKAmkOsZQ5/pKod06kW6Ktj/3R6BsBsIZqbVKZv4Srv+CNKMhfRaHJVPaKrg3F08MR6qKrv
LWItSfyhBp6z0526Xi0MI0QRWNlbGwz4MH0dxXjx4w2c5L5e0kHEnU1b6nBCd7MqRwLPqIqz4wif
uNZTU9k/4aOJPVnuo2BODVc8iDWIP8cCzCzoJOZRd/qPJT4a4IvSbvmyiBgRDt5AhdDnwbmSW5JP
wubmqGx9YF6/uNgqtWU3O6gqmEj+oEfNBK25Ovx/otoromALSSeajkRtWqvMsaCweYWl8H927hXE
/sCEFavTz/ONTJbSzqba2IAKjV1D3kHmTxU45oLU/ZRtC8RXH/f5v39Iz4Adr3K6CRu76QRjbTJo
xIiHiWmyNpg0h3pGsppOVKxt5uKBqbZ+t6ZwWXO7034J5mDsC5J/GD2E5mnme/NRiS89mY9sXjIg
87i22en7y4boniqTE/lNIwewapa3DB01eVzrTqp1GjpMr7bGU86Pw/GuRvqZekmM0augLN6bT9f/
16OLlfQJ1U8q2qPzar7EKudFzsMaVBv4Qjyz4nx2pZEbqGLCxy5geGST8zhtmFRnnzWET2iJSzsD
W4nR0dlscl1xJEj/EyMcz4ja5JA+87v93C38sZf9OE3Vgv13uiOuHXNhrUibWQ9vy8wPLk/p6/el
wYZwlmc++6OonGOOHx1EkgjG+d0fasHtS9lFPFWWy8jzKro3JpQgKNP6WSMyuRfOrJ4yV37q/tDg
ze8lph8gYHx6ibJFe+Aql7+nx5U0XOcdof4n/G7XZg+mgQ8KPq0XIpbhe6wkiCRBciRmyt19RFSn
aW5099rtb23j7RS9pPYNF0jn/4viz8ggMgT3D7w+XIIWg0CEqQxzYBdRhI5vrPOEpEx+/YDF2/ov
4YA2qlJ569rYq63xs4LiupVA0Kj/Bk6eZbMFZNU1NWhFGMUEXgKcI0waprle/CKm8JgelDxcD3A3
tACRHn3Vv8BflzXY8LPDb9cgjjoVjZfi+eXaAmwwc0YRXV8f3ZJYbfBPufeF3OooHqZrqMyZgRq7
8mS4+OfCoQT0SwTrYpLYdCXX1IulA/pDSlSzl39q3WIx2TqUw6MRL78WTOCXR7ssnOhpXlNcI4ON
imI+dnxnX/k3N/L0uimIFyLxmgRMkf2s7xf9DTE+vDmK355CcA2aP93dXGkCZDP8iZ66fjWKMCIC
tT51HZj1b5/5aNxtzxjHUqIynLQlafkDJ6GARPjXPMrf3PhQRqB2qVEDDJ5XyDK3SYmRpNXRmxms
UNPKE4JZw2/OLwhbPkq1uWh2smom0V5T5fRCSu18BS0uTYWM/ILamDeBCR55F9hIbWexju3kjqT4
pckfxvMO2oW/sFq3aki251B3dtu/y0fZBmYzUxi6lCuqhY+ws+Zigm+2Bynhq4roRWWOF1DnkN/6
WYn8OqyFAE7k2+vADppwkz3FRSed531LFEGiHo6B+N3SeMbJ4I0CJXWUb7tmEqLq8ih4SVX0wFsr
q+XPfJalU1Jo0OIkx0QSt15BNKmXhUUl8DlACOyw8B8AZ3MHiqvZjM93F8z92L17qY8x78HySnbp
GFX4PnVJVrVEETOM4Kl8MVktQeAgZb5wlb/kMtxBtJn8GtkTYvQzS06yEFqModxzxg+u6PKo1fK9
LzKlJBezBW14kfkG2hZNykhUN1TNGLEOTnCA7czpXb624N7kjb45ES6K2brIeqp6Dn/qhYgAdxY4
xj2WTCwxPeVfLzOYEEH7vT3/vKJUiPewueEbTDn+nltHBEg4pYQk/dosexF43iGQ7CWt0iZTOv1O
sdA11Zz7OYN/XuZwwRliix1dc5eNmifwaeDKMCR2tnuCk6WKQ4ahNA/lhmRpJLVi5CqkiK0mdWNV
BP8DA3mGHhENFBxJdBTmyCkRef1G2D2iPJIpIq5zsSCZkUa5BOj5+AzHn/mlAMikR4aC8HXjJNh6
3l98CtWCduVY1AJltWJxr17sIeOBiLkZKmNFnHdJa48/yn+2c04YwGaL1LoHdryyD88pMqJ8iiZw
Jw5m7KFRS3zUnwOEoYvTuRisoTCsRgEEm0cKKg9SiVHjPoT2zWKHW1wOOxywxYcR1SWfPYBdM0CT
wx6tb2Oq94hg4x9s0deSHJPBm0SHXkx3DDmwQ0I59zmQi07oc6XTUqKxfyapOkNrupnUP3vGNyHs
xdxMaaK/515AQU2All+AQKNVdoNfV4B2HrIzQ6BTLjX4dJPtt0hflV4KdaSqYtIQ8fhe48LgsDi8
6hWua2oh/9I/hxA72ieI5dSjMCaWT9/yuBSsEgFaqljr8979Q0qYiSSE+j1SrFwFAav/6XBOaVGZ
/T3WheR/V0pYlKHaa4NPBd4JrXd4t6p77ufBUByfSXQrEOr5htBYhajE2mXsWi3WsMWA+GkqfTZZ
EXjlzEFxKnJTaR1mNdl/Bc+kMfjuBJQBdsejkNdrcG570EJ5BtaVTPZjdTL5HVFO40ABr+q9Mret
0QnWcJO9fKKA/mYj+JQKiiezIjd4tXpsOOCciWblq4+UbD1Z/4gVjftlecdwgjpvwq8C/GJ5sR3p
2EpljFQbpJLofTPLL4TM65uWTEu0i09e6tQrd4qTPJcgjQAu+H0fS4TTiIa46//3oUAQYZxF0bwY
XoDBiGJCvfmDzg3xljk2RY5kHCYp5jeeXAUW6yPReHi2IGcmvbemOaHNsbk/uUsRGetiKw4hd447
svEsZx/NeGTNUbxXRMFME4duUmF07gdYj8vgLFod+az2SqybBB1qI2skI3Zd15B4HiLnSNmM84Sb
O9OylDkibH5fvEY+gpYnCvN1qIJzIUEyM5r+oRehcWcOgOV3UeOEt9qeIsLhjp5L4sxoLHZfZi25
klBXusgj7nwNwPRvHJoOVGMa/HqKT4497asde7f5NWp9vR5JgQWJCqYu/fz/0EI6mIufUoLoNZZt
6PJiX6+gRerAueedrL5ILWplV7Nup+8IM4Qove7NLt4SKvZG2/P8lnxjEALeG1geJhJzMZNrC4xn
vFgksgznyfe1ueJ2IKDv3NhoEcFPBtXeWLcYQWw3x0q/Ww8yZJytE+eOE16uyih7FWPQ6Tst1TF8
R80gp7ejWZUSaY69F2UKe9H9kFcg/CHAdLCLnxOe8yxRBROLZT/RPP8/IqgOnBHLSXIKrsdBni0b
SKnDvWPWOwClDkxQxudJOU0+H/DlV6UpuP00AvrSeaTtO6BEaL2qA6pK3jXzdIQZgNdXr4dx62Vj
yki9GZ31ryR0Qz7bJ36zMCjGgVanwy3b/HhPfvwCWxOF42bbbBPXYdjOUN4RX+PCbByx+YThpD3U
vEPnSsL2I3OGzJ3OhdAzy5/XFY1XbifkUjzlI6cktgYMDCjEib+28ggzx6GXENzdW3gj+cMXX4fN
Vt1UKLhK6rV9ft7SjoRYA8JsjBkgS0S5m9ZR1dIV4C0ugfVHys9YWrRiQ8xv6DhXb+l6f+YHGtxL
gQE/wRu8t1W8W+eTcV3c1sxf1UqmFDV+EsJr9FrCI4rrMlrDvhBxiDzJz+nVT0X+uL1p2PEBr09M
H0Fe1jdYjNroXZbH67gSMdkVi8lKZqr1yO+A1pN/FQlMh//gjl1WK3mRQwVKjxqi/tSy5rqCa9xz
YPNKhY5SFeO/lqlo2X6IJl/gHWtSm2OrQvk0UUrqxX2PNxTav4oRuIC6F9cDSww0bYa5QCDCLavP
LwOXVeOFRg1njcuunLdzpQlCjaFsYjYD5Vbs3dq9H518A0QydD1MLF1KYb7LhVw2SF2sjnv6kVLc
HWY8RTv+SgAEsc8V798B9NmOoBaXdePSxtHZH+Y9OU3gswy60d1tH1ZSfm0NbxeYDTdWw7yMd7Oa
0PIAImAAulAS0NGJH76wK8ZSAY4l1Fq27YgZiAzw1fVvs7+vvhSXsGviP3MkJbvzQE6txfKwhIrl
4xKmYpGOVSm5MXEez9EPzIN+o83bfaz6eGzTH7Z9WbX9gvh28FtxzOjRPReKpGOz/fcJ/m6VclXb
Pz0tCQ40q4P0tJt1bWYKTnYD8+LJrz0aSDq5NCYzEEa6I4wzaVl8WKHg1D7129ATr+fvhvoR6Ncm
EBjcnsWgJ6/MmheQiDSZLEzTj9vkxArYU6WV3ruWvLZCd2Zx4m9gezCTVlPBvuLRVkCzQ1DfMtHg
hLte1L7v/2PXYmYI/EoUat5+1jeDSi4ze9G/mb5lfVFXKlHuA4fWVwumkwgdAhE/ZZ67O8VIOYeX
uzVl7dGVn9tUYpBMNN8ELlyjjzWG5S4ehhQ2nCDtHZlb4ho52KRV1mCjpQxxgerbMqMhzwVw1pYL
xqwc47l/ogjL2kp6xbSU7B2ReKrfZ3FuAJJrFEXMEGyUvbNKF2I7AjJBtaNfVTCXKE6tdW0ZJi/o
mu7Sj+tBIXU5dlY8hvR49wRxGRhh5O7EjME273DOXex7qwl+Y94VN1q+1/fPK8GudM3dSt+V//v+
6mnmoFDQ0QwSdMRmLHCZZ/j2gLrdsIgF0H0CmOL0QGN3lzUKMVhW1uP1gfZmakXHTsZRxVlInk7f
QcS71N6NX2wg/P/FxNvTDoecUrLqCxeDdt5bjBGvsne5IvdoU0TLgyXl+5mkIrFMYijOYnPtaBFK
wPJLRUhHjxafzMUe3FmiFOfszZYeDhho9K6F7TN14FB84K1YUV4AqYDvaGV/WZlFguEXJX4+wVem
kYhPtZ6xJn9hYa9pJ088rea6MXgmmit1wHnnu/R/wUk/qWc+70QccjzR6AfvSKQ+h+pM/EdN00WQ
ujVjzEEmKRaWfgD6u8sdzyX2tQHtOYxnrfuXuQthMtx5vq6Pa/m4yNWmpuUj1Tnmoy6O7+tyapS1
Espp35za4WIV1rNc0aL8A4/chd4lUdDiwY3v9N7JnStO9m/LsC1RuPx9kuQRfbNyhuD+lpyt0h0T
XocvTrTxqxiBjDOVbYJ21j8bFMkkWQISzcTEsjo9ryCyNTOxpwK5/QrUEVGaX3DIReEp7uRBktD5
MFres5Vq8nNI/zWGtGUTCewz/a/3bpGCKiEdPpHfWdhv+xispmgvnZf7wnfnxldeyB5nv75g7tMe
vfxXnS5nWLaL2uualUr8YIZpqykltpANPKrZZmH39tlWQiTd45l3yMwrR1cceymm1a5f1AAmq8Nu
D3m/y9x5x5ZbB9hhTewlmbTl3P6KglzhAMS6kSqlayAu+f5BXTwaQp/pdxSnOwBs7hTtFxDFmlr8
foCisEyN7M3F/vRJXZpgJj3hrSSHqrqlYTi8D3CH7QbBHjp4lcS+7OtzU397TUSdpnMk+x94RMav
XdNSkxKSDDxXfcq/o1cdu54rh/ZxCn5wfIJE4ugOkvwsAQobXA0BQKwcbIc6kiYSh5bk8lzJgYXX
QixQoax0fTu+0ghVBiX1MGaQhyk0PimuF23f0NKip4IOHvPVKKWeu3IFchVciytNLJVtRmilFI7L
/a5Y+260DwCe7ZQF3HGbxFKXe1c7MALhDUFejBsNPlbEvUL1RuD2sgydRQJlKYKq5AXVVjqpqLl1
p4aruTOOEd28lNg4Bic9jD7FbLIitcTKVcUVCGL/br++JJ/j3z8aPWoipeRxPgQWOyhWW81HGZIB
9OA+PyyVu7/XAO9sIq1Ux0tAOh1/b88neVSnLbkztIvsE69quBxomCnX1RH8la6w7/Og0bZQHdyq
Csos/cAZfstc/NnYHq8xp2GIZX/Bof6zL5efSNWUFzElsSMq4rWnYRDn7cCTDVIUSjnX3JMNhdZH
TJk7zJIqcwuCCD/g1J8sSToJiRnXZE5NqIYaagYzEqxLe1jdBHnEvsL1tXs2gj1DU7xe9DodQy3u
UxHPLehu9xD1/8DZNucbOJ1wsoNss5T7qvik9FVABzb/aeIgUAcq8GkOU/NtWqzkotVPL5tJvjZP
Iq8Zy3vXt9Atu1FbfhHcsyqvnYmPSpx6dknmF0a7lfyjMq6OdOFyH5Kuu+WVDBNnH7+VSmFk2XHd
X01oVJUaIaAOxZ/qH9duAvw0r0BLII/dL4Yi6OdjagzjVitoiP9eCrWuUl1bTtZR902MMgw4n65J
cCOSfw0lY0vkhkW2zn+Vvd9XGmfC+thgkWVoQnvyDbPy85JYeQ+eUh7cto1zUrE2CQRcdn4A9axx
hPDuDBXKaDdjIiVmS7M+T0G6ODeoFW4oBmCuIUkcq3rbZbHW3maO+ynpcXYGjCsG1rGqGCRAlAk3
VHF33D+V4suPh4LiL8fG3C5dVyzeVtqeHG/F1yz+5oot4YG84jQ9Tut8pCkP74LEbSZgzVJCwTAx
RkPCAF2/6Dr8TaI5m6nBIJ+yeVg3ggVS4E99L6arr0YSIaWRIHPyWxIvnQj+FZZHGTifZBit8Sgv
EEskETynTYxFsM7EUovWo6f7XajvvSPHqcEwYe9/ZzAQZmWQ5OY2/yE5qzIFvRP3nri7Lj/lKqC5
v8ycsBjpN7vAtP9PVOmtY0hHEwS7mF8Xm2xeklSgdxjwimbyplUmWz2M+k+FmVnsSIe54i65OhQE
Tn7EPDBOcoOmWM2J6ZmUKxzmokGDpajXyezei0UBFp2z+viq7z13PThXe34fz2yWjf7fTWrQIumc
lcQg5r5jCGE0qy5P0XTP468b4oRG7JMK/AdWMtgXu2rIhJSJefek4xac1JBCaHzTptjEKRTyYnuL
Nh41Giq3FmsPlQNtJwEk2NMtfwqOmls6l5+nlWYSQ5rEpykrnUbkGTQyzvDUvnfR+FfV1IN6Ws2e
K+dZapc/UveG/NW1zulHoWUUJzKV4lOjWbcih+BWw55eBtr0dQpjJxHM9g9hmClOIfJPdvqWm0WL
W5yAI68TzsVXU2guBtjDUOWW43PpR6la2u4Py33HO2HlggMxBY/0ufA/shsKmhlPQJCifnb4KSe0
NjFMjhq9e6W0GjYweNQNlGudq33J6dRmTYsvNOkPd2QWGHWnRaFcgnOR2B7DaZqYZuqVcKQgtdVh
AKSuJjzDtD83a23qPv2wCdrXR7QdGYPZLVKddVMFF8+RNZlJkAAoNM7bXRU2+qcjaqP9RKxx15j/
xkmcwGbv6fnHNjHlywrsS6NP8QZzloJAxYxlp64PbJDZdIZdjG7jtkXbO5Hd7UpbFOL3gD8dAfb/
t/MTcWuE29z1V+ChrNjUnUAFT6GvtGOgbRnLcD0LuvxW/UkhdcQ+k4CB+ma4gCv75W/DdcxDA4WH
/jIa9CQ9oU8X/ezUUwfYCJ1pFe1/ZAr7dUSXz4AEYSlaXv6ZZp02emg/zD5gyIAF2b5IoHrb3vra
3AOj9EIDHqqggECedweg9KfhpEs/vi+qMOoShcNtqZeBEQsOblyo2aJv/CNBPOBvnXxb7YdgKIo8
fdq3Pz31O7pQXyCIV7fAWY+QgtzirJKfwdDkBj1pYjCFAcrkEY8s4qsbHfHMUD/e4/bMyjImlqWV
9CObo2Oum1pgf1aXUDg0oAlIN83MtBkbIOmgFWGDLb3kLvINDR8/AwvhKsnhA9QQ1+EDQ2eOwJiJ
VvbbQ9XyM3F/G67kkl80L17k6OQ4m5NM++4PThxzaUNmTN6HBe05YULhOMJPfCbzjiaFm7psl4y0
C2syUMbUqmzpT6VttJUKobaYtfK+u0xDeBFDwEKTqkE/j4eKEteRjSDCoJJjdt4n5rw2Cw98a6p0
zMGsf4xNekAaHcXjeQUpvPYOTknlJOLzVITLULUkbIKRDmcvPHFDPe0JaBVcgEWQu9apQWb112ku
JZbaPfsVMEpOFnJ6zObRp5L30PHasxioxlsokvLqkE28E0tF8a1bwY9eIWlHVrXEDvQhe0rBxjf/
IFr/Hy5v+UNjQnXOZHcNC6R3WFIUk4LYqIGidZjZYEKwKaB68OSug7mYKUjTmtYuaJEsBSsMUGwp
Q2bnARteKLtB/k4RYp6KXCHPcDSk52f2ZSTfLGRDK3SJyG0qByGi9IEH5GOfgwFQmZEtuhDJjAeQ
QVAqVea1ssu51oJx4zsSlq6a+eK4pmRzkJ51NDL/XFfophexRYQNJFsdACRpdndmCp6/CotJYiGb
Myc7nKtrSjMKMZ6XCavA2pQwMlKVNL4I6BD3yM2Db2v5ECq7XpbNvGPv/m2BaOW/LfzjqgstQT/Y
2ude4uNw9PjMbzuzrFqR+CfgxwGu0dZ6AYZfSaLD/6rGsc5PKgILOV4PiycjF0KYkHhzodOlAVA5
Z53yh4BMbB5Hze5CDATIWEVsGCJ0bZKrzn796JfUCqEnD76IQW4x8NVLGG3MAKLVEcU4b6o4+ScS
8ybgzLJaI+nJyeZoHM75YwYeM457E/U9nTcY2g4JnKAxjdK9L3t9PrjeNHtqPnFL9zHeWYwhUtUx
0BeO6dGTzWy0xxHj7ZShOP7KsqWqW7C8wnw8mvc1CMQXEDNVAhuSJqfXnJWEmhE8NrcoQDcePY1F
bSCyQoNOoLA65WO1HF5zyupjI+sBUA0tvgAO5xr28rPfpg2pML2IXKSkCF+5ZBoqgCvjaXZxmm+T
XfQZ+2cNZAWULkCHYVAhUXHvxQ4EknDsC0p2yqzquZtwMwC7EzlftumFtW44xc9cqUVSNG2mfbW2
xCm4PvcQQuZYPbA7upZVP1LOT6acAXOyXkf8bLE+4eZWEeY6EbjN2w0KuAiZlk8hFhqzNp2+JAnn
0ehKvMyTSffYG0HHFMvAmdkwl1AE7dwgBi1f7iijSmJChEJDUi6n0qoFNNEwCcjtGaH70n7LnBtY
AM/zIEJCLAkYUT+u8sEqY6GG4XjqOEIP6ujpypTdeEyXk710drEvszJqEnWvxr6SoTLzsJJErK0t
p9XLUdGpfJHGN0bzmZmFXBslFILpev2FgdZHgybyJIUzAV09XKpDHY0wh7OHLBiEk6kpjSpoKgdI
bgszOSBMga4+0CcZ3VvmJjRBUJV1lYqQ7sc8/VqVt1Y8iXPXzsfirt6+4KorQNYVXxv2UQKSRLuu
l6/Trm70g/d1YSENNisZ8GA2yZ85F5u2tX9J2GzAzJ1f+CTglZUkll/YsGwmbaWYAz+BPxBcCxE4
T4tDrwQ90yZ1KJSC/wy75n5UibxlLTr3TSSH3PJajQukXmZc4xMZ28VEIAuvDy4hUKo9ZB5D17Z1
UcODVVRh6wr4Ry4AvQFmMdc7PoXuk14Bd2Kiu1GnZUR6KHYc+m9SjRV9+0rkW/hm6zSmSoRQIOgN
C+3KJd6/r5k0NFXvReBH8gIAwbJg5evVpHxypz0tQBCedBNjtt8g7KLjEN9p/0nygL4O35+uhDUQ
R2CwvlBAJINbXOgWx4jWzIRyp5mpzWvMbWkaUq/80A2kf+oM+IzMeN6ZoMVqYu92QG/8W2MnF9lD
gFpX6oa7pEPkd/0IZpqEnOLAC4u3G+KgqZQouv3pT/iA3Evc3DMYvlkRNVCa0EPoitEttHYNsf22
r6Ztm6adIA4x5DOoxiTfaYjXsQrCc4Kd9wuPXngM5hMZhdTesaaxU8Zoqrf4ZVgg876NJDV5wnIV
1sQihXXvB7farSkFctdrMDihEzAEwUlB9EeJA+mQb7CDtXFXZIvL+iqTPjFfgH5/HXSTGQ4GEA8x
poqWQVjGQ9nqhVYFUj0ANIhdvezbSL3Um6d7asOFY3pb3dZ5G30rZAVrLoHpXtabbPgfZ8cQXBZO
eSXrUZiLmChnNMNlslUHSbAw9f692I4QtUzPbOd5/56A1pTSzQAbt7QjTG93Gq5DNNwdvUfWCTlz
GgGuClmEaLpGW+Onf7lpiifcUVaDQL44Zu+DoZFIA7kutiiI+Aik9g7ZX4DU+sS0HCJQNmkZ/iJ1
AarQiomkYFVtqCaFDJbO4HmG6q3Ol/9CIgP1f74Q20dx/JBSO3YApFj691+VBEYWIQeAXAslh/jk
XbOyutVFLGM+Zktzt574zTfowaMDIa9+50Cy2qVfxZHPb/WH5u67ikPmFLXBa/RPjSgE1taxKuVU
zi2tiKbYRiZCk9Jbj9Ya8qWPTgFBrZdbR0Byzaob7AWaZMbfOF2mB8fw5laa8WUyma/NM7nXiOwC
HDOMrLw1s0mYsFm1szohrv55Yu3pfb+bZnA8/KpLexOkgL2h5gVMXYoXPnnSLNEYv98Hg7Pz+bu8
VPOp22az82JesCntVYuj+bSz8IHFBUdt2EQBYs23SpDgCAaP+G2zY9jF3MX3FHlvT7m8ZdOEqS2h
wVlafTwqvhLCozgzOBUfCwDCPilPEELEq1QbczmjTNIZ3r50bFk1PtpX2SwgcX3DKa5zcjCrEvpi
HSE4x34eyjMi7gNT1zlYnMWFffmCfTd+reOzuartXqbN1uQNWBQGh2LlKIO3fucwhtWHDBHlYITs
9ns/5spa/Z9WR5EGgIKSxyCYOOkYK4BXUn8gzkQpZqzTSA97WFPliEa+/V5JjcKJD+8K7KY1MJdf
JNCqTW+t2w4+eXQrimdCmbrO82ug4v8pKawCeT1jP1l7PTpCeIEats1aTkqNkaXQq2x8imofdJRf
yeE9TPO68UPKLdRPiDoQmOzYQZjRuNzbeHfD5dYxQXwdaFlejW4sv7+aEsCcDX11SCXDITz/Uzld
q7MsmcWCON/XiP5QagyGUsEYD8HLB9LxirjkQCoEu2xBNXyXZpXXcNcwzF/tHwWU6tl/XcEhB5tC
+hnY51TSzU4EjRzCJyrI6fFWO91ReKdz01R1b+2Q2ygeVhGV+dSGcpD1IN4XLbwHLNkM/4CeZZQq
QNcmTkpx51tmvKLqbrNAM7bSCYWd6ZnKVHhrXITwi54Lx3RNzNDtby/3md3P9I+t/8kolWijH0UV
N7NkMg2xCKW0IO2BV2+YWTmcltal+o1VG2cIW/LfI7XlRh8vJGz3Qe8xEOaMKQ4vOJ+IJzkkmTj4
fa1WioL/JAQqGIIIijuf++TtPF51I0MeDFOmhHTsxj99PBgIZjKbDlj6TRnGBduo/9hPL+3r5gxl
KXbl4BeqNuqjyTHqt+pB4wg2lgOj+FopxA8mcKoVusErg8EUfAIpSrDZ1MOyM3fDcbIq48NQ3RJZ
44sm/HV5yFwxcPFmhoFdaVrjuP2VVSAcPim17jUVXZKguun2gYdZwxRA2W7+X21qCGpV87wTZr5q
JT988fNHJoJ1JFfVGM2mJl4KMFb8Lq/XbKya2TKMPfMXiHGRDcQWPQhahYmjjGiEBp3QRuvOmtGj
X94AqdzESgTQ6Do4ajmhdiNdJUGI3k/q/njChjnXqUDuA4sQeEMh5/k06ZGgM7/Idu/khuXaqCF3
l2Ltwimw9g1H4+GpUk7pDo6MCACLQcsexAoM6ymWeazlBj8E8HnbYVZMrBahYSG5OhYyTRDJzlK2
8OKIar0/X4T5aAfSFbgW8fUnZuwMJjnK7sD6ewY4S68sfOyLuejLhgaBbGh8YX7GWF4C5SrzaLVR
gCp1RaDrMXwYEpvWcmiLXSKPSyxIA+WcHoH8gfz54dq6FL31Y76QxpMStwu+/irEYSvVwJzgAmLF
p4mYti7yFOgzWno4evCF+7JtY4u1OBJ8Me1BvRQzHHcpN596Jsjw0hdt9KaPSFrR0uxXoJ+N0z7+
f7PK94B4apaxq9fGurbAEOTjGzHp7zbC3rnUvOb9mtuaQ7AMwR+e7gIrktvQ/KEmWW0wKmfMF9nd
H19FtHkbY+eSFDXcG7/j9zxSHFzWGR/0UZ6Xmw5uDfqb3qfWqwcfQzvmLtjL41nslrADGVhKA1GU
tHDFf/nL0wW7WHzfLnLP1+D34w4yWOQC8afjN/s7MEI/rOSrX4I5XTsRromaQkh6XUlIgg5ULz0E
Sa89vmdojmgK9t7944FPq+b/5NLhgkwC2qk9UpoU7WVkZMXRKx/4dRpc2sArisoODGSAhngdb+Ql
DD6MVaABG3scVZEjqaenkgK19Tqwo8TGuIDLv5EuZAxBIgLQ5KcdoBEMHn3lrRpj+AJJoo8uFz7+
p7bZU+ezvxNs2Ck6J8bMYBRQIP3w9uaWYl8Om0Cwv8R9Fu1Fvn0YcxHQUJkUKceYicxIVutnMUQp
WoIhsOLtZDizjoQo/9wW2HTu9nOOix2fnm/SLEsEYCEWKMHwa3Xi7o8v1s5oS34vx7ytfx0vS9ov
O2j9fSK6dIjJMXVs56F8yK83SCX9+aDVX07dSt1c/hKpL32JSKgzsLBfnXjwIBCP3fiNH3bTOTem
0O7K4F6PHdGoN8Lvh1UofNB3AYKO7MvhEiNLDknqzj1330lsxHiu6FNxXi11bDBYFIrVUALVHceB
bYpDPZzY44eOj5m0htHQvk9j3bqgBCdf6e8YAyrQ+qN3YH/rtz99qP2FONJwjgKAPQxUZDPLUdLx
AQt/JY3lnNRK//N0/Kbmgspg3b8lepRty+Hmj0wyH+tKSv1/yQiZ0T0ZIvutM/K55BVAsoQpI4mj
IqMNWHOJHgFE9Yhgt+/7zz53Wbzy1XBLW3POtP81Lnp0pd4Kfo96LTb+invb+jBqwUWzNAoigu49
VpVUvrbRoBeG/M39CEC6ujGFrYkDikDZnJc6adOLjw/RStrAk/rLZW/orZ8B5GdsrwZIaC/kpKy2
JtByXSePHOOyFFzSGVPqpChFEmX3vFWjeq6GhKbxK1t+47vPG/KZ8epi5LQAuiK145OLWDRWITXS
0yKb4ELLGF8Ryfti+TKJKHlaJhY7D64tzCXwBBR/zAmcsFWBcusnUbdJvGzJ2Pzdk3ogqoRfM27p
X9rfZbAhXJRqjXvFg6jkHstsdUB+uk7cYnZwsNpChsg99i7EXBzDyFquNe09gOXsOc15Ucf7ZKbP
R+78OzjhrdHXPgVJzjVisMCirfZiiFuRNzcm9iC3UHSzORTDn90dZX7IPus8WIfPksj7GhGwM9oE
APsYYq1ilRcyyvib9tInMTMx/t6aemcSypiYy5YByjWzcEZWykB9PimwqN5JavAIOSrqMBsMZiGi
VxDPhgWgaQXl9oR/u+0vt7UhGlfB/K6X8YMyI2k0m3v0y7hMZIxdzUd8DgkwXj5kh3EnCb9kPxrm
gHJmTWwFliYcMBadgjaV6aGnBRglwuOwpD8fb0vaYO6tC0ozZh0T7iGYA6/1r/vf3IC32eF/vI/3
ZNvicKe33P5hzYLzQ6PsOY4tiBvlXzYBOO0zUFG/IFONK3k/6ne2/DcwQyHaDyHEidW7DDtOzQGR
73Cx4+vnFr6h6jJcqolZfPD/bIIwCoUqd8ISA8Qcwb/Nw6D+Drz/eVUzg+ZULulBWOxCKc7a1+Zy
7sOmcablJ4bxsGdB/+GpkHyiolMvNyT7gJaW8eVybSd+KwRy7qiLqZtU0vbhKAKtY7LV7eeNJIIs
fPNabP5/QGCzqviTklN96bTsB0B5behc0dZR7ttRR0Y9c4CSYH6RdyNMnIPO+BGq/NCFMQAvQlFu
pb/5vnET29c56cKeJ4RNgalCue4NdWiuY9hxelGbrmZBFPTAkAdIo/KvUTwCwFf2ZxtYdcEivE8g
SAdH4AvQjiiJuHV/JIfswJdOVrz90BLnTBhKoSLFp8BIlVlbxh5WCO5UHlKs+KcBF9zs21eT+y/k
qcdcsRLbxxvuYJof/ttYLPWAcruzcZjGDip3dtLKpf/6MGEpAYNzNVxhZrHWfCcmLSyrN5L0uxQq
lyhE08UrogOTst0jl0jqBNZt+1ayi8zY8TxJSrFq0w4bLimYRBesbBHhFVljDyfTZhP9t/hOdMFf
TAxLBm2y9BMgpwkuixQdCAYg06dX+QNVNUarsOuFGYJV/8lpaBqQb8Ymw4SgMznFcUxnGRp5yUen
TZyuFMuwEKALTvhPha5/8XCIBWGir74XBJate/NdL8JYXiDaMmZbA/vmfZg+n3WeGi7XlfMR1WX1
B+J6Sr8WWnv1kJ9MjzTbGRkO3NLym46DSyiM+fPPSKk8F+askdkTADO72Bvqo+zIPyohOQ+2DvvT
JoZxA1Ce3Fe+NQPHC7smlZE4LoFx12b5ylVsXuCz6LYj6Zx4q7Ep4S+cSE4W+WBnbJHhEmKue7Sy
nI6N9gle4yIB4Uza4JU1EOs4mlm9Au/np7WXYDrqmFFvONMwmDfZSdnQ1CO8WlTxuPBBTMeiaHfa
y+19PjfViczW/dVojf63ok0RwvW2vEe2U7s7tATxVx7nx/aaPAqIQ3cZvV7NEvyMBiLyU1gA3GNv
FAZm/Wsw8imQyyPzPSyWLqzJQ7ktXPIQvlksaaPHgs/g5HhQTb+iA5FODElxydWYemUCVZ+g/SHK
AJnsUBwVR2M0Qjw3DifAXFK+8JtRSnw17JfiK4++nBwPme6GrlnDN9mTo19tXy1uzatLoWOBKtfK
9bAVNk1WDST4uCidliP8QZz2ikC3vIb20qgpc5KzEVXHAouj9rnuf6tU+gJ/guAS3h2vamDGL67o
DYeR6FToGp6j4DeszjuTMHDEQkURQ6PKpoXiClgiT15odIq6LSnWSNxD4aNYqtHQ8ZhY5FFZ9/IZ
ZnZKNg8ElaLjTG0Hn62eoOrqsEjl/YIhYC7W1PG8yvzEY9LBCxQRT2FBpXcKIMfspy2epqtQJtsN
0L/kel3k+o7PidqKkX9muTJGI0aVNjmsDhwtGfJkbYNLM2VlTtdn+f8v3bRjLpVokS1tgQR7BN1/
4+cSw8KPgnYMXlLVzTmE0ILXGI4RTbwMSgXeocQ/U7WWlGyuC033qUA2pojlVG0ifdVR/RIznaoG
u7m6OSdjhpRBnM7KyGhQRd4hvO5W93vfMHbH/K/Z0M3aYTMuCk7r8rgSYvoET8qFZ8fle3IEMnkv
lCSj5jTNJodKuVx/QoUC5NT3fDjSlUWVv6a93TAWUBDT9DK+KJzNGz8IB9uzU8NpoXs10znukUeH
n1tJKpC1+/f33La7dbyisa/wsz09OjQIwGfO/qzRcZT0WiGGEz2F6LTauMDEEePAWU00fjdLqCu4
scIPG5kh5QgnvHEGVPq/yVlqYvnvBZizell7RO0Ez+sLZYhH1wNT++9pXatwnz/gHPG3gv0AYPhj
CCAc2jj0bTN0uBaeq7DlIpgDO8was6aolxcleaOberqgBmcetjjaWA4y7Ei9c+g/jZb61xS3J6oy
EJc2M8wpberQxm/NCmsLpRFspT3YfFE2EpIEej8nnOtv9Vbo1xg9Jm2ic21VjeaqJoE2+CX80rx9
G89NHW5YezJDQ4/DY6Ka/rJ4NvzKHJ0RUGisBJNZSEReG+06E4Of3WMokc4bUdIoZPZhllprXbXi
rtnSUaxFTN4QX6jz6dsZSs7Djl9JtVagxCQFC+2pegJRpRMvxMntk+yiSR3d0DINvsbiM4cXeu18
Tqo++BF75xbY9LeCFcumtOhVNUVp34HAAFk6WNynMzhJz6bkyQrOUqIpLQ9o2JqiPx6jOY9bun3s
ipzHl1OICu3fp2vVou2rzZrOkvUtgsfVc8cjHtk7N6YiDC0jOYRrxJctP41dA5XSU2tRD0GU5+z0
0VKi6X3rRAWKcstAtzyWGvbjgNnPwM2xGhVf8ssQHISInKKBboSZ3bt6vkDTEAPnQYj6FlwuN+On
IxtVuZcUGD6QGkz6foUgI/26gaOlSmTZ+SVSL2Ywu2YMDYRcZQhduMWly2PkdwvqTIkdf32zqR0u
6e3McjayClMTdWOn+IfSS500EYWHO5kIj45ls+C+UEshzT8aRGWV+ph2JzimaQ3fHERHy5yEd7mz
TSmGmiM8IF0SoFPDyofUwzalV7RsjaF9l/Q8B25uMbdEmbihhoZUoKZDffJRVOrMGHZ71geOYPsq
toXs0KoSOs1Sblb9eX4+vo5zk4Efo7x8nWsHkOUzfdejDvL32v658QthCLDj5pmBSeMF+PIGmwVk
P5PEQVAXOimVtBbXtA1D2eSRDDmQTLdA4PUhhHYjIKtjPewStA3v3i8RI3chMKH4EmxL6CJHNOFA
qQbqpfuMAsM5fnJ8ZAdcouC+rDL4gwrh3pBdBdeCkrNhAd9r4xHXxlQZ8Xf0R84rV+V5Wh+LjUuK
Hmg3fN0Wf08qriG5M0wvABz0rNeSNN2PndJWxYLpWhsFoWVjpavDop2c7YwLrNWVI4LTj0BC4/Ec
dF1qd9sWuQ7VwP2GSqOa3SzGFcy+lNmkMSmf48RnXxp4foGvIB8r0LcryGucw4/E3GPrlvWGek7X
ErzDdSCd/XuaxAxtyMpqxwqcMMd90XvGVuSGbadp+bLQdpWI6OlQ+5kecolmdQbT3qjqf4kB28BD
AwmWH/omU1vRDaWmqTpqBe7PpwhLEAX7s1i9tiUtUZuuZjz4EkxFMWdRvENcEMx/M2NrpcKPAnUm
4u194ldbH/kdK3szUiMCIFjso/dihu7UxJKBq3BPsv2JpfVSOyDXwzdAQuU6cNztUDQTCyxQnx88
soO++JZ8+u4Qgcm2+D1Jfe3c5s+wKrrOQXRp46Nz9fj7SDyLezpRqV7eeXnY44iaz2I+ABUQzNw/
hqEAv97PQHVDf7W371yn8/l/+IE6m5pSQdabgnQVNN+BMrbRgBW3CEtTYd0hvlyyP29PPJK5Ucfe
1NQZyIpGjxCaEMQgeIViokuzqmXpp7KoRDmCmTJVguFp3y4QEqZTSzgEH9y13dK1G8s81SQf4HFP
7/6LM04VDbvXjQpIPzlNDuiXIG9ALoYjP3OgOCaUqDn9WeuMsrXXcfsyc+9AaSgJQjTRyUKYv6qI
anfKIKU8jwquP4zV6h5ACg/BE4uXzdJfs9PSgcWOGqZo7IZ8rOKLJ4rdvvIeQ68i9C3MN5kG4aY4
8jy2uiHwWEd2Z4sLkhph1uhA1yEQeOWGlX5MfrsdS41U8kAF9/nE9SoY5tCloJTWORwqY1xWSS9f
o8CUZChMmwSC95IFl5Ibav9b8AnvRkwerjQV/ZckmPKP28lnpAVoL39jTpsRmI11oTY9YjILp1wg
5YJfJgtgKgM0pm6GnZNRjG7igXqAlvhUjtMvJMOFS7mlIdJHOaU8MBPox8y0BJPCLmAZ43ALEaXZ
1e8DnatWBsykSmNDt13lGiy7SW1yYW6VFOkmi1ZFtQWIN2fP9Can2kcdjJdNAAvfAumB3Tpw57sH
gZoLcP/792aj2An1qfvD266Gvv4rlA6ar+IkYb2Tax7v/1B2cLCc65BiP/ZI9VY/VV6yK7mhaB2e
NKfMEq88zFJL/ytlOJi8bqxoA9s2b31vdJYHBITnb9HQ7XL+vCOO5ggM934etobsXN8V2Kd8Ff5o
hgiQAtNVzjscSmIpETx45VNgioTBJoXIkIjZuhvZzoAGws0xHmXeEeGlxTWrXBbFyRw9HOqY3mTw
f+jD1CtyrVv5SvY7IAZC52sSuzk5nFfxL7bQwr7VnTi5zqwqUso8+KamgzHCLhAx3ueVGxJ8Db2A
HdJzeplrI3qyG77PmmB0FWJ2ZZHikdaKzVBKjrBsz8hsTGssinJ4PHkxZfZA8n0wslBNqHYakXD3
Qut9yrDVqAymNbFTbehgCXjAFhYuAcQkemhDgpMuOTyGdI4V18PeAi0QbiFrKNboewo+cVJTBci4
0ZoHiv/Fzotq/jw91FtuqP4ZLOY37mXsqXyYcE2n2Hqzq2yUVJavCGQN2Id4Cq4pWy97NOwpiPd2
Y3oziHKx0vqSWiS3oo37ML/WY9rVzdJU5LEiDlZaAQuKHLwASjK5M8d/n0DImlGXe/grHimrw/ve
yj09xAIM2kpSaG9kjIqjNqlXwe5hkr1eDzUSXHq2BGbNg7S/poI6r+3dReCsPTNJfQJVQXweF1Cc
IGXrhQww6VKhFm8TCe/HrJZiFwOzVswSRU2h0IgJ4UOpwrWqxw88kPM0ifL4n5VTrjhdoZrue/cM
uZ8VTXJJu8NEMn8Ms3nVPS71AL7cfcxmOxhVHEup46fHRcyH1Zm5ei4hOKZvpaIAuuoaGfSigjCr
Mh6/MA5DGCMTCHQxJea9OuCGJDdPqo9m9Yf3dqlFCRqhr1MEXFh/AaLmGQsGU+euopnx1CDnms+3
eRkyuKI+G1MTzY3V/3C+h7FQQG/zxbiYyXiFHPayZJq79/iTcYZh0/gT5t3JswcMseihFqupZS+8
RaXrQeV/dO6rBdSQCDJEUMI8Fh3T/y3iy8g/cXPu4eLbP/5IQ5Z1nRZyl7bK2Y20zPVlFDekDh42
vnCpJeF5+jqDCe+MjCI2pe0q9KiNoolXLb1L+a+is8WwBBGD8oooxPxkGZubAvb1TciVSM5YKl0U
+p5u74lQcmw3fSOCozoEJWzlxThf05emABQMj+LGpO+Ik1K5L2mkbhZSo1CmO5sdYxJjsx7Dc7Se
hsHpa0ZUgvNSSlHq9RqX0iWHg24sJpoR85uyNp23MYk0Ibq5oxWCaxrT9YkCnCJ/htyMw8M/ntNS
bhfxYKvaUa1/u23zwLWVWZOQiUOA0oEbvgkiexjf3SNRxy8fqtYEwjKHAJdoZITcgBCUXDXWwSzA
KBgChqA8mRZk34U4zQczzWtmWMRZJRH86B9IAelOfDEVddpy6t70u7xdnBbnn6PqVQOxo/oXmPjz
1EecOu04aUk10FPwJK7MXoHaMlbYkXTY7qoiEWtlG2QQMQ16cjtpkWVPQlc70mb2e6oms3qBw+9B
qklYukz1IMGsP3tpd2anAChG5jj6BhsKFnE0qb53/6KkTTfr7yX45pGvRX+AUOnWmjVwO9FvPEWW
t3F36sAFTSAmtLE4l5FXT36g/AaMinbrifphXohYKjLucD7bJHc2/RrSourRGvCutqiSamn4wDpj
xwFAtJqqdktxS25cU4Hyx1OVrxr2kWtvZiGO3ijp73MCYXTMdBi7SCwPHge635xRo4PrGTOpMNGP
nP3W5zSVAdMarLtMEFnN82yLskWj1LXZh3ac+SkINjdXxgCnJMO/oXJjm1dkJu3npCtlmMIlMDid
2sOwqKkRDWjbshXf3Zm2vy3R1eZkc5n4TgMAGn3GNekuyy8afSIHC4JvJP4eVhqUakUR2x+85Prz
6CxSYt4Kdx9i944y+CyNVzZmEX0fLFYqPgGdPrQOzp3JaY9X1174UGHAlVAMfWuxhR/tkST9GrCf
LyoMjB8IKaGlVZQDOxMxduvuOmNcdVxHkhCSfPbdRUR8aa9ZRP9oeXrSEVYPjscIhW7mpi42vIQs
zUNM+VC5kjfBfLjfaMNNQKgupeUzYiQ0fon58l0y7Izub6q5qBZ4ocNaxUS1Eux4BrITi3Hcv4Wu
1MzVSJueTORf3vtWx/5IVGYznb7fM8BiV8QzP9ARmwlzelddIRpedUr+IGLplZDVF4VPBQ8PTICd
7xx+AGmMZPgLusWzlqJnEgVRbSRrfyNSvYQdugNHxE7mdgTnWpq443+PZ7UqE7wuOX84iLo51t9n
Qb8Vo9fi8eUIw7BRljagxkDy2wFJyRXF7+445nGouYLtE9fAr0Qhc/S/ngw2zwi5JiefuWsKlasZ
laA66WUaSGukIg/4Sa+d8+bju5U8/o+CJEdxbV+/Zv83XjWcnPVgtTbVtr86LeztU4rTABs6SlkU
uReHhWjDyl4BGT3X3FX90/+PE+mEPV7kxiyA0POIIYrUbmU6Cjqxi0IUueFLrXCcpUula5IRS65e
yMrNuLti1UmRecJONfjZ9GJbTEv50tUkl8nCnHvTVDHVCGu1bAmmMwNeH/Kxdrz1cEmUyWIUNrr/
DEnXJDNTv0i6qJBqk/OmaIc83ZJGCs7iLr8zWfXWFWZqL/gN2i9y9JO7Wq5g6FGo3TFjrR+2t8N+
MUCQXyKcd4VbU5xnagCj2Vy0h1g6PfQRb4v6pIToJBaUs1ZYZpCexEu0Ue/WRIt2qZFbtLW2dQyZ
IwqfnYg9569YquDkX+U2nE1II0DJB48SobwiXKv4n7X1BRfROiuddWL9i1SaDrOHXac/3xNLMOim
BHq2ZLY0yfKCt95r6LZ3Vu6S5p/iINImVWBQ9btUSQtZWaXIIwInafTclchPZHKXBFr1WpUE0qsd
bHgvUUzPqOAijHq21oc/o4HA3BHGptlUHzQNWazKrrAENHvObYW8cOUJNLPPm8RLIFJHlZZrT6Ww
LryFjWUZ7hiDE92MYL/WK/ODCSyliRf7YhzaSD7TGijalp1kfcUeLJ580dHnrpzYf3EHHg7nk0hl
uVcVk+ek9nW8PnaLQaIlBj7Bg3I6ggNGrAJTJd+s9nzmLUxFFIwjkRfJil4tErtnhPULJt2hx+Kc
BbbKVnCEfDk9468qdKX4q/LVOkUIxgyxvZ+hpdS4OpAaWSQlwzbe9ImrmEOgC176NqyHeJZCXR8f
rOueNqggcVsfNKdRlksOg3CdpRQBwMvRGW2gnvuti0bg4UTn7LVZr1ELD335sPQtAzihEE9wESyc
ThBxIVAoitPN2PgJp1AT1nG1K/gcnMK9FCR2VDfZE2Vwk7KaKXUp9Qn/dD9vVld/QF/6dSR6ZjHD
p0kH6VnM8vTBwSwS5DwOTPMvYgI8U8iX0HEHb4c+Po2Y8NdPsgMoFo4Jc0cqN+GFrz1hH3hzXg9/
O7He2yoT9BLm/BbgnNVWiou7vN7k1IHsPhq7vFLvM4ArJ+74GMulKjvOhmo2yWPKcP6wyhfELMSS
pe2eF3j5qiTVIVdgS1hIVc1Lzza1MwkcO68WYtyL64qMHZcpORHhcM/cTOI5tDy2ptecU0nS66w+
4Ru3e14lahyp6Y5xdzoRYjXbiawd+1NuC3122TYV7ZL+D2qlDur/Pjnvq8m07jHQxRuuW+fcbTfy
iNJF+OZbpTw5swbUoHzSR/gOKFgeJixnZzheLhxgo8iGHmzP/32v/CkEBhWwOpmPUK+znAaHtIDY
Acaqxo+5Kzit2An+6d0qRI5UN3FEXVSX3BYF9Voz34husLPCiRgM+n0YjtCOHWAZ6GiUaWiam/Ky
Z73cX5iBd2bpZDfTzSEHKw1yhJVy94mvtpIfgvHwFCUBq6ObHB0MyZJH4W4NVvliVJdyUn4O8bS1
o4bdxmoF0YMtDIS+ewccAgkA/2VEDLTqV+d4JHNPGQGZqK1ZvG8TPwqgT6GhCvRZ7SxeyepBiIiv
FpdWnnbfREdkJZ5LotrWue5qsYXm6qSp7+rpewTbCLfacVz65zmwG4u2dutpf6k2pGVJgquqrxfO
GSAv/9HNf5bxZHxHwKZurWKWHbGkUbUOhR9ieGeztcgreLhMR5ipIhN8CCVcDEfSzJTW8SAGw/Kg
nw65srh1rC53DK+HCr13sSz/WLAKnWtniGmgRHj7vbMMDLEuGasZiPWTn8582WOkjQr9G5kVboHw
UtL32pXqozfl/To2eAsWrVj6RaE0ZSdrGvSZgoQPbjhrT2wM8VSkqn06LwoTu+bwLdCkGwfkf5+k
1lV38pVoshLro43tN1wBDdLSnJmdw0V0Ux3T/fSHvTy+rr5/TvoKayVtBtLl4VVNweNm5NoteThn
tWe7Xg3v1OugWfAFvcZTUo6A0Lpo0g2OPEhTcbvl+cpVhNr1yAUBS8ZqDcyi5As+1Ik9fluJ6Ka+
6izD4QCZ2FMRTGoG/pnToCXycjuh6Op5r8DQ5PMtBSrTXsULwOAb+jUUY6FLe1R97i/XyUalicCy
o7kN5Bb95nyvJxtr+H5Chikyjihz9ZqpL9liWh1JqvH06vvxwzItwW5KHOliZphUO4y8YqAZLU0H
LuCMoZMD8+AXOMgCTihMEDlAyKQHg9Hj/ZozjSFRSgkaOLcYli7OHpuQf6N/o43Ma75mmqtACcUT
eVdlGGmyefC5yk8lSc8lTYTYxWyww0fuD8h1ecfia1gA/48eu1eRrx4jEzDL3zETMKO9v8lKuWAo
Ko6OZqHAybK7BWoqvJ4pR9Ui0iVqIRMvT57anqYXpzj/5S2fflBD0EE9+IO0h8/5VyTp4t3NjD+a
RNvw5Mpj4QU0f3uaQxDSOTd3ghiej1sTK/M5XZd7AOKH3NDySFQUF5OaKbuT1LcD5vz7NxIwW5+7
4eVqKoplydNJqRZHLhCSoUb70SMaCS5LHjW7i3xmh5MurMQ7HZJBSzBWRfQA/zEb0MjpH6k5DmUT
bC9Py9OE/EMDwLsRHPQlDIFTP/GjNBaq5x2IPEZalK2mTIfDSBTypdB3OJIqFKUGwBqFvavVQadA
TdhLbpBLXuaaAE1JPSNfTTDWyD6LEH+rdrIZH7LCOmHD3fL0k2LS2Wb7CbBbp6L+RSbiYEOrJqGh
sAJhLBccXoxhvsBShcI2WvYRjSf5w7KKgbgqnDsTQD9Y9+qMn0asH1wNrTmoNriCNr5L/i+apLdP
b5nbQKlSu7mBSLU8kOruZNovG39zOGkySUw3o6P1IFF7vcF22PyiMIYUlEgVWVx+CxwY9RbYn84t
MxbbvBejRiPo8hG/HRztOjEC9a0kf3I4g/KN0lGe3c3z9o/cWZMSrnjIr8hn6K6wOe6F6Y7ND+3p
+2S0DKAfBdbCxJ7vvFZK8rBin6V8OEhNRfO9gUJdp5RqKkD762x3hIUF3zAeSTa08NU3mAPBTAh/
vy2aPaiEWzwBX79InQCD1Qu3RL+yaGZL+ECofNyYgE0RBrd6hyZzXjifv+X/l+dH4vyWKxiEbwpE
+Rl4azO1A/CbRG04VReTFVrSJq3pegOIubBf1PSQIeT+kaV44ic3UTcvXQBd791I3WBVBgvnTANn
0Y3jf5Ef+G1jdeMzjRgLLkh3J97rul7d7cz8dDUVmByqh7n7HNzDhwA2Q085JE8crrCJjLyxFfXj
pl1CVrnqYvu3IIeQQ4eIk+ayFY3RaDkbw9vBQ7gID5jaTIGhpb9wFYSsSjYCIlPmxQhO4mfFGlIw
Vg8u5ugzQWwhJHF3LUY44CtDHxLcY8CVaJe9EfMNHrJRD7ROcesTIlFNujRA3Uk+rczuIGShrWOa
qwSjHv5l2lp4whlVTOcxrOynJHNcCZLfr/jEdufcwKeEbbsr1zOTfHTotLwh5fUNVx4hnLTHzJzh
wOZPiVgV69SEKOS5/HVAB2PgFa7KFEq4r5CmhRVelSj9oew4o6xU4phSH1M0E4WNAzuONfe5N8jN
yfFn6PgEzHznM45/TidU55ez39AWHIR1MkZ38S0FbXYb1oosAzHZpffR4Oph/ufogI8xJXEIXAxm
n/KjWtJg0v59DWbdqTVjQ+Jkl8FCcRke0vDgPQA0ZkTkdSCqXv6fTskqEInD1l9b99AmOomJMb7R
O3wqLwUNsCBXNST54gwM0om7rpQnWfQs0HHW9MlqkcS8hl+gcAeqoti9KeEWXwkYXEPoFPGRh+TM
gZmePbsKmA8XgubwsoifRWW418nkAtWYz9TmyHVNW+tvNmIip/e0WAPI0KEPcz2R6H9nERydrGuW
9R/BlK7+08dS43678lka7GM4MWyny0WTGIWz89r/LwULgw/SSJcPaGHQcPCmR5spXt7+or96GHWc
Tc1baINBTA3ymblE/uIZh5WsQniXVf0NC91kKkFicuOYYCHc4QdcNjeTsBc2Coo3Fl1w/tUG0o0S
FVZntjMIW/fv4f1vswrOvasWu8o2pvEcidTIs+YyqejN/lBf/i+l62eKbpE+LXqmFyXKhauADqRs
gGwnyvKHy2kovXiHOyE2TLrqe7H6W/YZImJmM7jGuJdf5SInnAEYfVmd2Kg2pm4zEZbsKurOkF5F
fBZZDKIrmIsj7XncS0toXc927RnYRbeAaQDZyKL82rd1Ht8QXmS3KCxErAhJuaC4fWd9gqWH2Neo
1MfS42yQ7Zr/o3POXhSkznsIDgSPwUfn9cdwzptfM/5Tt8mzgHi64sAPtyFjRI0pjC3yUJ/JYUII
6WCauPpxcElnsQZs+BVuk3WSnW78fl065Cf4WEqyTCxBTmaEyqdbOB2MP6yLs+GDHEULOoBL1UOg
b8aaWOnnyaaoJpQRljyEHgPePgLqVuj+SN6dZgpmdLI7UxIP2imlCyjOHkyBj3taP8lYD7LaEu/B
MYZlct3QxkMegYMFj7RI0vj/1zluH9VOtSSGENxpPTVk+GWBAaKz5xcg4TaOnkXXbWYLdXj2Bx6r
bU+m1PXMApkf44LPKDNysg1dDuFohEN3R6AjeMnrqpNKVuJ2olQWgpQfkc3y7i5D9Tk8KAJ1nFpF
HrnoAn6Ygz5DPSjkYI8H2PQMib+wujhjusiMX2CX0xmt34NZFDafKxj2tBxZjDZ3rot3iuyNfYPD
eZgmFXi2RoTeCKs+ADt2sCacSFGmv5t1Ds2k91jrOs4wwWSQfBePxRh984wCOdTm2Md5SnKmTSIr
xu9r2i7c2WVWepwUMJoTsBiJeGUA8o52JSb2ELEnXbTzilOMFMVtmbyUwDHHD4OfN6RDxC4byatS
/SP0bKvegPCMk6YdZaVH8VWZL6np/EVvnRDTZJdVXy9q3DLe7w906lBmwNhF9AVAk4YO3tIADznJ
kZ65U4Cu2Saj9bmngYT+CMg5FrxOuWR40PSsnC5/Ajzcrms+5iPsO1xm4GpSXXU/twl9AKWztcoK
Tzd5ycczfpKBTSRvXeVTtbRRypFiVNK4rsD26xR3EPef8q45cyEajt2a8BX0TJbynWpHvtK01uto
fHLOq2QV1kji6U+ezAeSpD+0wvh48LpPzExQnfkCXSz3+vnDtQPm4gDo8wLjTAx+yuKbVV1I33oW
e2afdTdQmfS6iid3eOHJebtO9FRdiQ4Bh4zudgRT4NpI6v0LbQiuUkAfQ5P8tYR1hUAO+Daac3yu
HSBjTuOg856/Pb6mO90+jr+AQwYgfhfmSkYq+Z/K3d30q5OYQVG0geTAoDB21UYiWr4lJDzDiZwV
ErpDZlNzyiXNUASyPTPNodazDReQCKM8px11Fn12vvsZG2A+xypPZUiWW83SEzxkMQzqkCIjjhhl
8w2otzAQr7/YIzj2aQgfB6wzSvGq6c1PlzhIqNn5oOBqpxFEw7fUM+1CvDMQSR0O9qaI9357y4zq
X1LvvsAu9WLuZCehixI4M01qNZWSqfYZ9LJhmzxXIPi0zq2JJPYXI66HLlowdLrv0fCjh4hWKiRc
KoHpuEZD7WP4g3lC0YbT0OdlEkx3Z5y+FFZ3w/fupMgsKnJ60cUMBIR1I2DBaW5mk95/71moYpNf
uNp5BLpe7q0EP06tFhF8otuaGrPP6wySNltVhpbJL+IO6ecJZnKoZbj27peXwuAabgyTYLwJM0IB
YRyW0ba0WdD4CtHjWUdZpT/6IVQ3yF1JaELK3T/uylpp6g1GyI+ju5dhFIVX+7PGjiftK8LGlgqU
fW2TGJz6rwbQ80926kmRrmYWXL2DFkU9fyw6ZEVF8LMHAUQ6g/HrCUrf64Gob82CIM9EVmljukAF
Kn+GBT/CQeY45QHaUCBzhQFRpEV9+TqSqbwYnOB/XG5F6AQM/sGtRVLLF00ReBsS03Kbo7Iqmi24
c8n4l7RCFMx5i55vYrWKzd++3IrjJho3LZSnqEJWdWs39zSJgCTU9CamhSQgEBNhIAOYuIIFZFkW
SeTWELs6svei1Jzb57Ntd8fnyC2UINcH3U1xImS/u1+m6zj6R63QHFygcqRSSHquGSL8M3SRbnop
HcPGW+8C9Er0Toek1yCNUAzWyZLciOwU2voiTqV8bSER4ocNZar12U2AVKkXS2wwqjSVXEYCKM4J
bOeZ4ahkUV45U3/T1YyXSwcS6eWGAyFznPFa0yNk1MC/FJCfaL+bHv/tjtvlGRB4y4duJA5CnuXd
4PayGA5rLwbM+A2eHTkY3cxqTpv4oMkBQmlXLDJ9BJWBGMaelCYZPFVMpK4U7jTaEyW6UQo83UoF
eLMvBePYW7KVVqa1abFNGBZXH/5iOvgNl1oMJ4dF+NyRwXhnfIw6yxLOw/qVoKz/MTL2ERUv/V02
75kcBAi7K9doCkoCimQVBV9voZcuQYDqF6I4NWmSAn3sDrEJhtMMt65Bm7lQD9Dg9cRYv0xz9Yx2
R3genbsI9OkEcCnh5JlZR1w3B52KB7agZwT9WY1mfJmk24lbg4HDcd80kbaNDJqT/mWuJJuriIX/
2F51BmhoU/305M+72Gib8ul77E8M2YGKUqq06yNZEs0CLNmjtvEprKHPqvauPwpGsTvehWXevQ1W
7pbJAVEgorl58vKiELNvNMVbKbSdmgqxG3m8m9CbHJZAAhx4sktiYO7qBGMenR2Wv/n6SqKE8WRd
VB9jke4Ec7ItZ2tH5VXb/zHcw8h6oZFmLUwfSId6SEpY96udH+/VlDHKc1CZOms5ThTkmTYQ49Bw
wkQvzZXSOrzZ6rq66agZM40w9sRm64CsOfhwxNPGruK3jftUlRy8rivg4PcEx/W3lFpVYSoB3bkv
3C/4bBCnLVJ49hoPW5i5JY7EKMSsLoCYP+KQhEbmXpl/UeuH65zu4P5xDCVrRyYgyGL37VQNYgTo
0rKrXJ6KACuR379aBvqKRg1dqPa4oQ/64gzoGuR6OJb8303vuBWuV79nQ2Z+E2P9SN5zp5uMKNIN
LetR1ISRV/4pIqKinPAJpeBaT2iR10LtcZtduJU9arMydoQE6XMVvucTNgd/69LGEXBbL8qvZulq
u6Ql/cmsFlU7wCDvl2Ou/V+KhIxRzggR0o9idDA7FHnsKjmLXRy8ea17lnNWSC7FpurAKQZyUCh0
fHjBN2Dscqn5CnbGJ6iQv+11Bz7U4+BQMtsBsl2sOFuIY8LvCcFo22nqvK+uFy+gdZfUPVRAsxxF
MUh7Xu0HaIg1pX1USaVGBGIoQNsFg92e67+jJ9y48P3Xp7+cLdOgRZfXFlBsnLt/xJ3+yiD7Ughe
dgfCrO0XUCbIhrnfMx/9tk8hRMUQarZZfKKOQonbncGtjG9Jl2T/cUJ5y45ySj5nv3LdG/Zf/ATc
g+z0UiWqeAlXWP+slbQIB2Zinwso+m8QfC96g9La0875HJx5AvoDP7pyjuzKr88mlhCXVX2qaBYh
x3UjJyX2x+d4V3h4B+NlTkh3pGej03iUhchjawwy81K1TUMZAzfxgY6gHxn9q+ZFFIXe6Y4oyJ/C
OLPw8kf7cKZ6ViyqidEBvIXNkls0cLj82Wn+xQAdEKEIig8bmlZhX/M1+3b3W80ORk9eCcvRHkV1
XvhhE04szURtx/IpQQJe+/o/CuayR76jikxKLjWD6SdC4SsUeeeMRkGHgIOICLXsQ+ne6/4ccEkz
r06eQt+gzmqAH1f908k0AaPh2t5eiW362iZGBU8klfx+Q413CXjhI/0/XQInvDrAapZQ1WOOoYac
AmNlVXieP9SLAWij8qcNENEm3erl+7Eg83SLoUtkMpWqyLXdFK1K6pzf4LD4muVSURWfvv+TR8kI
k4+yr53d4deKo2VMruwRZZy6xCrdujh3j0lJF/J5AZIr1QNtvfYqdU0UC1dscXvYZ9Ff5cUgtIIX
X/jsmXzqSqEnmBy4X9y7ugDTUfz3aBJMqKFSphx67FVoO+lC8MBz66HXalwvQbotzL8PdqXmmzpf
s9RpMs+PzJRSFwwb3Lx4Jal8ALue7pQ5PcmmcsFVI6BE8FczrMjPwWrRWTCKe2/KSurv653WUuDP
0DWstE63YodZeexwHisyb1Nlroh1C0GHmMg+fIaYqUmjyVZv/MCMSnVLttMM6oFehSFD3YxSOa8q
30QKv/qMnvaEn+feyjQJv/BRHTb7BMVvW811ZwtpDEBHnc/joYXTBaMuRfiLG0ge/oXrCJSrvMRm
Od2jaM1ygWP0+2I7zx1+rg73zokGGZhxglSikeUpC1RgvxHpbrbc5kAjzX1Yz7tBWDReWp9DkJ1f
pv45vDUF5AmZoSwC1Z+DxGGJGRaAt8wuZQ8kMWyxfsvzIbL2gSZG97cpmsdB0LhJxQjBzmMhCren
nCI2oKPKg/4Xfilw2vQBBwyEh0YWsmcL013sRoA8Zqi8ws2tXQgVXoxDcBI5A/AJu0qAmjFmPG6g
1yjKIpfHcnHBXAe5YCyVLBgn0bxnW1fNwRInURH8HUNtZDriupOHuNGmLmaBmlvN9dn12MqP6spJ
D90quv53Ygz7c+eDiBIYreddKHbkN64qOvXVInUy+/IC72fp+GU2RUr7u2oo1PJmZzvnI/AXv+IO
ykveXsl0xcG3L/pm8te1Fc/OoGnN8hm96BFoOr9TQ2WAccIP8m4EkmTa/n0nMmfqQM+JPdW8uNlI
54Ef5BuFpoSk06eF7I5VBaCLRwYADCvNJ9qyGA8wkCP0y7DoOATUA2+ZLo4kK3HAR703uisb3gFQ
GyiU/bLhTv0ogkmLC+wRoIyhmOZKKwtah2dFIA/YdwaRMP9tHprlGg5cg0R3wm/bIjbMjMyZf8gL
ObKYL63sPnlknUevi7jqFNe96dj2E16FoCiGZ3x/QyFry4Uqynl0gC5otUsZ8unnruZZg+bkvKb5
3DH3o2jTAf4F4SIjWpoZDB0GGeh5cuuBylTEpTcpLeNDXx+lJd49K2hu9ZOMNxidk8rt21GQe19O
n3A9MB88vtID1KXg3JB7uR6TaCAVLeBfeW6Cx+bR5ahk0CK4JhsRaOOcplzmQZvCTT523ynf2Ggn
0vcCm5yuyY1A8HAI4WBJU6OS+qUq+Np7gmUdYllCW7vQMhyG6f3Qe9H7zQyrelqM492t0/pixfZ5
YKJ6zbFe7/e3zYjEPVxDogK2reGEHXLdIojUVwf+UIEfzh4OmUBJQT9qnbN5cyQVA6QhhIpPorb7
eqLdPXDJlLezDLn0U54zR1CY5OqaL0kmPtW+fbLHxfIUhzHCkitvI6kRLu7tfvuEpcGAHTcLu2QH
w9jCDK3j3vgK/WZzqndVRQTZFZBasRcEpaF1257WSZURpzvDrw3M94DCybb+kBBub2UcFlK4QBQS
emnHPtJPjNixLtco5+MD5BBJxwW9/WMXPnMuAQRrS1dduQmYJRMiAs2ivslKIr8PGm2ccf5940J0
kS1vzSwgAfLk7XGIEPKUxE2UblNTrNXHD69VQAtQ3pnINxhF6Ao87cixZSmhlANgWIqbrIdXJseB
Jy7nafJ4bfGzlhFlEWcKVG3Byhj5FEPG+GrF/0pZjlFJF9cYcFZs01wgaTGcsRQjkG5KsfuXeNvO
kPTk9gPQhnYGTDQ51DOrAWZjt038dfM2t+NKpKZEM9asS5JY0tDl192+/yP3AhV2kz9ItB0xRakE
pPS10jwIHOVPjx1Rg7oLxFjDeWgrf7UWlGFMGTHnb9JuXP4lt7HNRyiZzHkuB1f45agTR9CFNh6R
h0u79rP5nN+LQEthBK2ec4TyW0ArfEOApsNwE0KA831WHwdNnquR7oAfnyE3Y6d3FHf+0Y77sLrA
cnxUdEtQKiHFWSyE1ixLA9WerycfSmq8C6cgnI7cg8RrjHqKWOHlJI5/loc0wSC6VKTuFEvPxz/A
Slg3iNNAkYYGKZBSqPCkM1QeJEA2yyMreGv6P/qsNl8f0jyGxUaApkEfI3Z2wfmo6u9xovVxoLGQ
rfGeqfKpSfGm+4vEbRdev6VZfr/EEA7MWYBUNqQOPW1gPU2qDBrAEQX6aJqqz/vIaptSOULh6wod
NAc+dd2NpfAv6mr3uoTTbFC+M88HnofwOoMBjnyNZBY3M+xWHTiHGsJ6KJcv6Dps0sk4Jf1zhTkS
BccnFaXKkFkFXlkITn0c0ZV4QGmw5adF0uI3NRnWkOQpr/DNGm7AD4YogXmNT4d5P1mZU1O1om7c
ctL7yat8kijOdz8FQYZBPzr+qdKVd4stN16mrP9GvJFtozgzqCz0w3WcgKKFbjS3h49vGf6G6Uzn
Mwt1uNBTeXRJeWSWe4zjGW8ZNM9+vI+gtkRflzPNqUB+OgNvlePStIQqTi72oO21TQKvTHNMp7Fx
NTqa6kpfLXevJP/Y06XXB1+7FkxvK0F/ZL7zYjX+FtNIPgR9WQhzuRgAQV0XNeJuRqDvnHsgDK4H
RR9wOKEPVtzB1lkalwjsjeo0FZbxqFrhLL6v2xYcOUcD8oDOmrFr3U2rgtjSHyZL+DrRKBStrOJb
xn1ooMm8/vVKV0rjVwi72cZ1sAve27M/dKA+o7vEumTqfM/6Tkh9/Dfkn1/cPcoyfCvkUyyvk9i5
D95d5yxdYLbITzu3HJWNU5g4lY3tLOpqZE1gbVHtKWy5abxtE4uCi8r1E+s6Nt7e9rsumSf7VVdX
Tnl3io2xJ7/vJNhfOIhIAVfpALw8fs8nLlXW9AEhT4eftL7hdbECWGutZU7Bn2H1u9M8R7ExC8nh
a/zuD5uOMp2RUgj9CWegOcnxYiwfDn/u7T87q96ifk52S5P6CxlZRJniGoqn1Ld40wPfHnQnIqrl
2Miau7/0h651n5Hx7gwEeWn340tIQmqSgUhLcF4YIyAR6Oh+XOX+AJGV2Am+c1bYIhw+PJNhMS29
7TaCst/r4O73Drsc/a/H8XuwUxwfq7c5gJr/6ismbIldlfjyi1QiZZGbpQKE848M+f/ucTpblBuz
o/KC3wBhdpqo46zUscaDuBG2q+4fCym3k5qynLsIMgAZK1mjqOeCoBpI9V1FGEYWhDp6pscJ0CiS
jpZbvPXhLRiPtqh5DgyOd8C+/qmUepB+540hlp6MYtZMhxTUYnvCsC0QC5XN/FkxQ3KTbwNl2/d8
yNP57RYj6LGW6mkS0fdCi1PtjqDBm6TgDgTfnnsDP8WzrJItW4Iw59uMBV7yJTl4SUqd/LKgyeNR
soqOKnuZ5+fQa8m2Y/tAdrl74+Jv993OMSJPioVyst6dFzxXT/PjYmgyEw1YQWA6qnGWtYTJxobf
9kl4YPiBzf4GOPIhR9oLLrXvvp8onWIg4M45Jrq/e/0jLOi+xwhwqjYzsasX70MzC7DIkAA4pTvu
ezWrCjUOZ4AryNo1N1Q1AKpP9zDY+KlF40gfbC0j/U0iU37CiMRF0CaaofpIEJdCPh/Jvv3sBWjP
KzZ4ikVaJuGS2B32tTuci3rGpKWOs5IBvfaAYhZUYoai5Q5OkpxfhDi4zz2IG6RiqFLd3ASpq7Fw
TRAmf/plwWUWOTHWRxLeKJAV7vto6tI57jSUEALU+WpZ2KCo3DYDbQKdcuZSD2Y+ZkNvRBUSV0pb
EA/CM5c1ehwhY56iIPc9OUmctwAdbVLHYHQZtE9ukRnA+DUKwVA8ojhum/J8Fs0aBbCLEswzav7S
BMy9RuH7uK4w6nFLZuRsRuOdNfXcI967dcVer0/gJkA1+E7zcVWdyi0YeWCUCpjVaCm+9DHnzMSr
DT0FRruUX61gfXqhg4lKWlDdPZoH8F8/RolmymNfVlfBLcnztfW1oR2/Z0bgYHru8tmxLBMmyglx
1XnTPYWYoV6Dc2SNuGfCftq6Tij3zTpeE9O68bOl0Az/BYzOkQ4QOLYoQ8cuJsTRG6/8Zu2qvLV6
5kjVUHl7cdoz/RxjfHuBcZmbT/4O6X2h3p0cYW7X57I3GJZN+vFNZkSRY6MhDpm4RCzFvi+hSJ5e
fJccLlQkO6cXLmPpO3VZADtDgJRPzZLsI/47DxIm9y+r/r1ujjrdrle3f7/Gp8PfHQfqcLPQowL4
bp6or1HPOBvnFU51UEJ3UsxxIKGh1PUBeJ0M2I9VEUG/o806eDPb9AOlbDIN35BazbXrHXZoKzUL
u5qgH1Kb4QQAjcwPyM+iP+7z8Y2Ikd2fVDe0N1cPLJ1CSDsIOxh3V6947WiSncCaeicP92Ag69te
Jqjeo1ooimNBMuK6ZMC8d4RyErnURlI9jJxZKAVcZRnXxIWR81E+fuHM9hyON9Q2NSZjS4buc0Z5
IPg4fPKLgawYeBBugsh8DIgJnLcDtOykkEnGFJOBLUAvZ3lf5UzcbPumvUvD4vOJQAIE8lOLmlP/
eSiNwN8ouluPNRmB+befigbSuidgxt/tUGVmN2IaDeYfFQStzRr1/GwSBmt5r/NxSNpl/H7n2ou9
gKXMJ1JR38JY8nYfdsjQ/41XDjWlfqICxmBHI4ONig7dZItf7irU3Kqsd3obhGT0oJewIUr2A+f3
sEFlc71VQT11GcrxFQ6jwqlQNQM0iCkJPA5TVqmHRUuk8D3//B8ZewODMZnmrtolz29fqb3OX9wg
tS78bH+/jAKE/kU1bQx3M8kjrWqEnTHvTz9fksJN/OWh7K4AbGklBLNLdCs4lOBxuMupF7PxQYJS
tZMQVudRpeHU25A7sQlF9WZsjebh/6tgKQdCvnodVJe60DSJcsQCP9GRqK7qPgcNvd4yjGMjaLlD
mbr7oLTj3CWTsBGtnaqZIhGP+zeJZDCaJfBSrtZT1p5aOGVh0EJJK8a4jBYPRrL+JuDCY+kS2zFf
qCg/LL94COK5xcT1PHui88HZdxSZDciHZTgwvPplkV0RwwGzTe6RscoHSf6ljaeOGfR4deAqUvBC
31Z3aIzVHotGah675iRMeqnKZmYcNF6A3tT7YoK+2Ktnr6PFEoX2JacJUu7ZsLQALAsyqaQkgPRZ
/CimXpVJN61dIRB92tBKWv9pzm0L32kc7uMkqJxNyaLR45y1NBnyjjtrUpUdsLZNYsrO0pfNohb0
Rd5P92gS0dX4Na8EUsZzLsxYeOHlIki3VQNrDKhaOC7dnpV6Kykj0Ag6sasd4RneSx0YjZnp6C+q
2cl3hRAfGTd5o40pf7/AfQIYGfomkzuM9cPNHz8OuFwDqvRG50ui0v7iX7jHIOpljFNV3u3LGN9r
dsesx7CNOItRgqG6K1No4td1UxLcFXN9nFunFR+Qm3jhhYJyWzRv9qbdxl5/anoBFUT1zuYIcY99
BmNYBuFlE1Y0lXe9afWqIzT4bMoP3SlDD/6s06A7McnnMtVYLwkoI/aEYUMiUygio5JwzcvfSHBD
w5/zVM9l9w6Qkk6PtN3g0d6snSad5PeLs59TAuDhGRj8es8PCcR34F2jaRcsHkDh/l5EFflz+S2f
QF96jNGE6N3wv4KwcRa8y4gzPojZQXn6T2PqcgXKK+XQg/RZQPRmVb6ayCqeiVRgsCfDMakWRANd
GlI4DcMWNd1+fyozyKDOtSoQmVybiE6mDwOE9UPDzt47nqFFtRgdIWWbGixA0gDOL8U8iNHKgIMy
S6FSqEofG5WRukcjgy1xYZvdjCD4H9nw1UcrbIQgm/kG1uC9etcuMymNrVJATdhoOXfIOB+g94mv
3A+3Pk7ypkjD42ENnZA1aqWNZ7a6CsF1IArWN75bEGM+qFTZgN19YMn9vf0qm7mW/1/ifA7nwTZl
Mxk6MxWgUfpkN9uRXoh+SRTXZ9Oq5p+BriTFVhl2S7Xp0tCVpjSj+pvrOTHaDb3RaqBkPiKjdtko
RdwU2eKifiUAFGI30qf3/UWGfQKzW4cihy/367H1IXcwJVkEsqLAPbcTm6KqnadwWSNr9p460D4Q
cNte2kW5dzGVt6dj9b/S5Tii8tsG0TSbWDmny4h7TA+AwQAM9e6wEQTUm+B9Hb1dCUhmY4T9UmCL
loqlIR4TnB/I1xiSJtVquYImTWL1XQ3OzYjdIjd4n8+qnYY1SXa0kqoopk1JwlgRBx+5vfRTID0I
nDILpmmuYY8KMMYjur1ikfq5nXKNSXAXVlYDk5ppZY1mkHdmn5usAOXxQpuEjZw13ggvZ9JJvgi/
mzx9bjD1zR53zfPiGVUXOkmpvPT3ikCuCHvRW09vQFIvqocWezztexMN6pvkHXPSbP3EhHD5wE91
kYlSzprG4zT0usB44rmUBxeIgcK5lfRa2jolUfhmL6Vt32FoRYrykbtW2AZNopII1Ff130LKH+u1
jLVgLz5DTbQ4DW3pOn0jsHLj32JMSHBrr3mU3cDWjgvUmm8SQ9WimjaeZ77D6+8Kr4f0POItgLu5
MyGoDMGB/Lw0bFIgrdWYrM8ikiwUr1G/hBgvP850pmnZe8pQnZCiGHxDZiC4WBNQhGcm+8zCaioC
ZDj/Blv77ID8ERjXIDpAaWXdht48aJq212LUP5aHG70oWm0QIY78o1Wkoa4SBYK+wihxRRFRy7bU
iGiXrMHLSl/dIufonU61X72bhxq+JjQukRZEQJ4LS5Uybfm4OhGAsgL+fQ7AObnjveZMr4NfSBfn
UgeKoen84R2e2Sr0lwu08WoU7GZ0AcR+VTzfVBb5LQ18mBvCEiIEHn9otlJFn3Vf0UbfiA8RHRb4
e1q3QSt7EuTWWP2gal08jNheD4RA9BjkM9dN552Ol4O2wjII8qCDYjNrQp3evU5mrUcXdmJUUOoE
8Gm4lxyaE252Vo18UCOykmHlDfpJ5IA3LiSKH8zU0N9hS2Gj0HYQ0KXueo90yLqIwUI7fFGEaMcU
c1+Fs+/tO5l6QZi6/oFlgdc3oKkkLgkCnaklvpsC1WotgK//3EimdvluPF63tTgib1SshoW239JV
3GTZJRIFYFqO5sL7v0ztw7N/yxUmcqxuhD1OnZ92Bzm/gOFuqLIFGff7v/TW5jCKV641ZcJ0hWqX
tT8Dea5tOWPA6Kai3hSDSMecsYFb/pUrsYxtBToJA+qrl/PPUkTiCfEmeYI7roQzZIy6nj4H4fHL
pVx3FRfxOwlKvYK/yNduw35YATmmwIlj400+hRWrQeCqaxkgHiTQUr6MA/nm6Rdhbr51A5kBSJSt
eR+eQJ/SKp+BCF6tV4dhfw+tAjEJWdXDlyMEQ5L719nL1w9FRvBsWFC8nRYGXiCE7q508qfeVsmm
zCZus9s/9uwndbSMhy/lbI5uT8/QKjHHjRkcqG0a44Xb0gIOJLPvGHzstL7VI5eZwq0Je5qwTxt7
uZgg2AboYsOK1qPgXPKdzm2sX5J5fVBRAORYd1O7bHqRhybMMz/xgVC7gqIieYZIFvF7qaE6jv+r
a23UQFNRwlzZDjmb06+muhd8F1NCLygw0QO5XRj7dIDbVxlTyppBwNSbdNszJzFycB5s6Dy4MpP1
02T0ONX/ihGuZwp8AbwYFKVSO3xv/r+lpsIubCruftxSj8pKqPIV9yCNhrR5v8oi4qzKDoL4qXAU
IEJaeROvKX0z7Z3bhT/tnS/a7/atSVvPJ2Kv7AEE4sSr5M4wqnu3Gw8AUex/Pq+VTafzMJ6dvJQR
4RtFmBOo0bsba8fuckMV65zeBGsAwPtKkGDgCsRwHWCSGXz1RSJeN75otK+bHHGDOcBLkqqCNhaC
+BI62m9AyMVyHpQbFRIcTC7jckRVGFJY8kTGMX4PYzRdw+tR/ED038gV1Amh4ckDPaTN7RT4BhCy
Rv2hwr4IRnPucRpLevXKytFwg/ov13riEI8WyC+Q4hxlaXCynuREZn6B5aTD8lq2QP7L5N6i/KfU
z5V1CEgt65ygQMwKr6yectAPGMSkCsCdcLfNaiea2eZm5zAhZFEiDhkkqYbgevUhqE2eBAIMIR26
Aceqd3GeHay42BZ9STd39Vq4VdCIYmfBSyfHSVow6XJ1IDxOj9K9EJF3wxsVgA+LFZJE/guU1kww
Jy/RisIW0u+1T/nv3ckCW/n6O0rA/dlziIzApuyOYxRGpBivCFaCZTSLMC4ZEGvo7YQJnY480BCA
16jdX9ofOKU7SAW0N7Z6MGu4MnBS0NzHmZQRYW5ubXj/R4AP7i4ZCVgafjp0U28kf1owkD/VINbx
eU3qYoQ0IBIIYjp39iTsK1zgCIfxVnze4UMnlRzUyZ2t5pxt2AgEyqRTjad5HmGLgPAMj3p7w6LA
TH6aD1dQFKdUGxP0HuB2jjdjZZfyWnCvyXNeMLC/bxwB+S+gzdUwft+zxdNU5WLa2EZ8t6RKwKaH
OjvNBWWFHjGE6n7rbl9FFvrTyuFZzBEU6WpNRGywLOb+K50XHy/9CsYKHJCJVKvqLnc+DGlV3ra9
jvv02B3wl4EeC7sXLUYksXx+6SEXlc3PiQK8bp07MzdQsIVfKQNYkUiwQScfsfEXngoysjVVf4Pp
MaPjpRSrwMwYYexyYZFkSmvdtdDfB6wg/2mncOhw2JmKN+9+0mRfF1jlgzfsR8cDkmxiFXWvkb34
VWFx7AMNXNnJY+6SnVz5b0r6UrEmwyxqm8E53NefqO41JgoExdFx1BkutcIgddR4wGLs2RkJHfBq
/CCdnZMFgeaideORrCyGEgcS45Exxzgd/8DkE4rczJs/F0H1m83WrsK6/DqHvrc1NYxaktBbwiOR
J/EHnNpqgv6cKe+PBg+7FT00czg4AOZKOQUAzD4HvspOhID9C0Y6vjtH9whgl8SbV6qYiXKfGEML
oJrMQd1H3zjPyLd1QdNb8REl8L3Koa2L6FqA7Qi2yeR9AXwLOafVpOlshKnvoHWynospEfXeOzJZ
2SW37SO76nFCmEGsyJQiwGXtiKR/v4BiVO1ovPRadPRSCcxZ5R+kVkRFymB3c1L/m9pq+N16ctaR
byR2EZ9RXwxMpvbxs4ScTTZZ1EjqeqSw1GW+oqR1iDrCbhKRS16v7lx96QrVrAIYjMLV7fPn2wPi
kNlSo4P0IFxIGMRHm9EJcJupsKpcG6mXK/PsyiufRn/HA8Pmrg6c8db9gDxamaezIR1D+brX8PcY
CHruRLMGEVUr2KhXdWAjyyz0tYXDWfTi/rdpQhd/E9CVYfp+a3YVuIzb+lAkbPv4m9qBPrXMKMxJ
nKJTWEL2upLf2ShzZ23atB4NhohwMtZXXm2ZmlJB3e26rEwPvXneDGUNVWPyw1BsB1yhtB3xJUvZ
9u4nSqf5CBNxlFqDBhoMci1jb/4H9D9lRKYifY+K75HIBJv7XWJdFjkvWPBwkOEKIHOTtIY3Alo7
nNR8xP/skRpzwXCx2QC+QwOOTfuQMKJc4f7xjEcmWuplY7dGiwqs/2NguT7nLsxr/1drbI4SFQnd
+biJt2U0MSY3wqv4bQILhtwmsj0dEZ/WoukUarsAeqFG7dZcNWHmpwER5KqLauDgvoS64gD65gr6
bwH/WEoKcP+BKTuW4Y0Y61thNJIt90wllO3kI3sGD1UxABg4YsA9kiQQUWRVzZ3utDAhmtAnKvqA
jpa9FXg7NcVflaZRrose7rpufz2U6yHpI6Hk94dsvdf7tiJ/hEDT+1PpMGEBTk4RC25MAKMgII3v
2i7E74LMGpCan0TtsyN0+jtBNM8lek2IugmqssX9++ZDZ86YgCDQp0qtgIaPIFqM1B7tOtwhWge2
8fL3sJSQXTdA84an7alzWsKWLzJpnnRvSsqkdYBkOLftJgWXI/yuS38PsajCDL28WQH0oiJsI8Gc
9CqfH4DZBJrI0Gl2pQc32ZN2XBgYvM0bI3W74p5yojqg0fn23Qf/svtcYb4whMbKvDEtY7h9aT6R
FJVZdoMExKCUWQ0bzxJNS0sQJb+2+onRna/VqjdcxmlSumfurTQrRlFtDcK5x+d2UwHEp9wqJT+r
LXr7BAHaNz3b0+9duk4/TLnzZajk4Da6EOeXXBuP3sBcqVDdFPuqmaV/uIjHHXF+4An5GPZdM41h
gaU+bwINcouvqy46brTKQta8cwa9DEYhDyg4nuYrkPkp8ULhXNLXRWctDS2tjaVik5YUH+TlrfVd
gUQ7PnvomkcH7i23HlkECBJEZn4qrGJBJRzHecpoTz1BN5nXRtSZH6XGnhC+j76Gk9OyI1jUPvwC
Tp79SAeaXqHfE/KZfwIbcx5ctgFZjwojO7ieYE1cTRx1t389PzAP0z1UvPsPnpazhCcqFLferA7B
jmetfVrUUOCO1KHa9kWtLwXisR+WZ0R0A+XdQp9FwvTQppXYmvbvLlAtx6ExrcZf8wZdk2ZBvPHb
kbMwDLlDpfawmiwTKqutkVvYPtPzsl6ElPF5Uc9VYQzov6YWQNkjfzyJq6nTQc5tZqqk/28NEjCC
k6qgCDRDhNe/GvKgPw6d5drX2SuAE2jmdHD2vhz6EJKqcYDJJ9vQn6VnRVI2xs7xbLV0YcT7tVJ+
KocJTO9quNWwrb7JJuAOrhUyUQXOLo6LiYoYchbdgsLjorafhgV0Q5C9BhjTebedWzvoHmUQIe+/
VhYdxDzllvTph5/2RXZZpyIZZ8TfHr1mjIdq0HBnycanb0EUoLZvGGf2+Io2dSL2AxHloMmcnJPS
jiz/ZhZFT1Fqdy87a87JHFB9QmldYlrXnJCec4wLhDDGDW1N4S0bCBs/ecVsTP5AFFvKLeCKT0CT
Q6oPIwJ4FUw5f+5vEt0KZTTaThLZ7x+SVMcqaRiQlK22Uimw1cNr8DiH7ATagdTztPz+o/j2POz4
AEq8Mi3q/podDtFjeAUrV4r9MTf44IiEhOxNGRLU5rNrN/Hi0jN5KZhcIPllzUScbULMNA2B68TJ
22CgTkCaQa8hpghjPmCWS0YLj9R6rWg59rk4ZiJftSRLv4hUTPVAEnfcDwuiWH9e78dW1fKEVITL
xu4JOdcE3X4AFMc6Oohqt1tFzdG70C/MR8A0b/j3Ox9Xm5pbpq6X46y0YQqr8Y8Tdp6iCfVIjHWp
QHN/PQVJf5oQMbXyr6YPJTkxO8i48WyALpGxDgvx8DgZ/QsOUa0YMEI7phJoeulzqVJmqZhqBcE7
umyTTMJqeaoamvnl3hN9zQCjzEg3aTrf9qDMgIcvxWJqFvFVKd3tFHSF7tsYVfIksyBW3bwWsIQ3
D6pmltoBWFZtwoYNH97UFjLp4xwpUQgRBgl8hBmizIy7ANeFiflTqq81lMoipF7NZjfNHOD9ST5/
cp282SdiYGEgUOXngcpmEpjWH8oemfH2Ys66ab9FJw3/VAUq6lPmRlctKhRxb+m4WGt4orOwgKTc
Qnc5mAB2b3J5IMoROQ2BrKZi1zAkA1p9YySeoFv+R6zfUTsyF1uy3IlmUeGyNabDtVQBMYyM69fN
mLtLBolUKipTPV9GccokuwRuCjDWHhb0NSIaFqtvQFe2CzfEY5UGhPteuDpUxM/sA3qhn6Y4rfyV
KFQv8A5XFt+fmKPzUDrPrdSq3lrL+0kyxv4olBBJeWqwfI3QPSwe43m2xrRb98lVInnfvFWqTYPC
7mFe4enjCVB79FtUBAgh5uRNGfIdTnGWZwITSG4jDBxjVhMvtkD07lEPh5fG6yw7uWY3lIiwYa/V
tism1XZxMFNqvqI2fz0BD3IQagJYb5rCBFIJCSoiEJjl/yC2NY2GlhPm3IKXsTBwjy7AqCvzmTga
Em2LTurmxht/+jqo+Ez0KTNiVdvKihyEiTtUPLm4aRXYtmSDhjOKCRPg4WZnu6nvbLcye0mWngY7
6MEGvpiZKmn+Qzy9ZzONvJhE09bGJtsaVpPFCKlgcsHpYcjNIsjzHB47oa95WXR/yL2XaWABN7ne
EtBwtI1Etr6hI1YU4AxUMQIlDMYdWVuWAdfqLJgn5D03tmK6QvODFWPoHDU4dcd3LPHc9u+DZHFs
z5R1O2ZC7RqEJs7d1HEybO5Em1G05xblxFg+76zYdEE0em8zCeEbTp2AxI7whwJ6Nzhpf3hOGmJU
xkdNcRe7HQ96Vm/4iERTthx68xRCuzwLR69c+/17ZK/mRv821hEnIqKNbsYRvYeJ+Rek54YgCblJ
7CCHhr43avzpH2qkJS6X7zt4neNq0+RWYoVT0SkZ2jADNI3DFemuUoWLbbXXzVdDqpAYv4saqzV/
+UUz29M5+oDZXDl8CWMR502k47OzxkDy6/Kamcdmn1O9Gtw5Vu/uARRsrdMdwawfRrV5hKEw2Rj9
cDEeGFyvEFJmMiTWjPtF03eAtFRQOUCtlMKagV+ozKJnKIOBEzZMwlbUIvllH5uUY6dUFhBBbxoa
iXkbE4/GWXM0f2Kgc1BnYgmnfd04MSBdsmecgqUCww2tgrMW5Jn3buVL5Zmom0BL8wXRwV/1vnmJ
sNz3wXUwUNvtbeXosiuFTUnrDVJCXxVkPCPai++rVVypON67xri4amfj9CO47jOPWsefnnWWgx9s
hVAPlC4nmXJgKwWj63xxgI9rFlMD22gT8ZitQAe43LKlYOFyMHhV+aUoVIFApn3T0N8fnVdKTXqO
xjaEaNPI49s+kTELVB6MGk1oAaFzQbB7bsMAibjRQxtt5xUV0nDZvwdpZ8GXm5QCiCRqPGHK1KeN
lgc6newyEo6qYWVX8scI7JGEg0G/zycie4ZZTcmtMQGXm3Y6LGKJ+eZeWeypjbLoS4lgBXeIBtKm
qaHIE2kn6Gy/1CWJ9wBwBqimLR4wu6iiNwLw0brEaujQlhssXV7+tir+mnCJQfNNb6njYvHJ6NQI
HKg80szkcHzK6gzQblS3fGIfpiRigv9KvdKHWuV4WSDYtT6RXDyQp9HcYmakR7rXnPw2bW2vQI9s
o7RKiOAItcZCpMZF5GEcet/ml1TLHpmYUAi3MniFbAnsRJZNEiBguCNgpymX/l8ovettYctzopFX
VjMwZbMAFp0PX7D1Z2WK3l19mJ0CRkNGwRJPuX96W2xddhgzghtPKkt0ZmiomoxL2Az81WCujB8E
K+5cHQa158qwC0QnWH49jQpV7b2IDMbkKdZEeIpFfkm+le662cjkjvHdM5w59PeAh4aCPhCliL+e
6ELOeUD/yJwmaujzs6jw+DA4YxxkY4OSoMFmC+ZtYR+fe/YA9zHQiznLdCWxEwFc4VzT6LjWPDol
fOyLc7jOMCe+T0uF6+6Wt9D8//oTxuh7YOYNWYK9iT+IRrlc/zwn7xqwNNzZEZASyxWHHjvB8vgF
PiN/8ppACiacURzF5aGz9xvdeiXwHjxvcLAM3IjCWr+Q8Jtty9gxNLnvB+QDrhWoEE/yGjGLsWjs
moGRXavqHYdGb7SaYW42YWztI2qGzc8Ll7c1lGg+aJk9p1R475byXGufan7pY/0OfmRMYH4HWpwj
ehXVaX0Z7l+/q953Bn7JLs2YUYMf6j7MSsUuVUwziyfR2AfG9wrFp33N4N3hQ7s1ZVx/YOVvfnuH
FySnu4UnZckfkeHnQopCdx+jo9u/fuXllWHeDDAC96RZVbVy3s+UkoGBuT6k20XTUw3WUI4tjrH0
Xbbh7oWfQ2fVjJJAZzL5qLHv0OtGVEXyGPDn4r9Y6dHtcHz/sC+axI8N28AjmozmYOzzvzrQLW6Q
ZDlVEuYSWlikujF6ZLHiQBvGLfQeYL7LMEr2ykiSu4BQx8nRFTQ674q7dQCB1xg+v9/xPEAKwoo+
a1G0l2e+IS8yjqYyJRzYTT8reTGGo/1LmMf4LHx+gutZZt2MzL16rhdd8fCJRAEGT8wXqd/q2R1d
mwZtY0308thqiqg8qtPON8MyS8Gm+Fx+SICLuJevSNc9x9cx5nTMFQ3q6x+7575zF5HEgH88ex5Y
ZBdkXgDRjH1S54pvsSKexW5ql6liaTtt/EeyN9y5JD8bgbHC8BqG6c2ihRf9F1Nwsp8jr+Tepswr
B991YSxefpkawyb+kcifgr5iIgxYHO/mQe/M0IPG9Tygdb31tn0BV6PMCCmEpS6xMiXIus7CNXeU
Gac4Zs+JamtRVWQFMpChwg2Jm/LqMQ2IWgkdOuStL7qoqZddm33Uv7anZtRAboWwv6y4rO9ySnuP
bu2+8QXu4gKXIXZXpQracV/Mu/oSUZv9URyQFx7BKwNNFzRSyZXS+y1uwUAJIU78aPoVvVM6S3mF
hciKCBGsoOeoXmD/wreyIjpgp3ZaY3NYSrOLH/oKIWaWIq/gf6fuSEvdA32YDRYen4zjn/x23TEr
2VRV5GOKUy84i89p1ASkRhiUugQUdvbuLxusAGh5bjLHPEQOSFCF4dKOT34yLI9JmMYq7iqNekym
X0wRE0T+yEytrBAHqv1UHOF5qrw5fDRMN7z9kF03zlvBBQAT060FZZ3k3NcGmMvqDzb4OuVI5ipM
imv9m6JevDmDu+MB8oVDgUQ4i34Ls2SIbmNR9QdLqTx4HGUcVjUaxvsB8SWXpX/WWztkQjla3//u
kaF2MZIHppzxFeh6wpyk8zOjU9N+j5qavvHCXMirbn3FyhkMFsU81HMqfY93919CiGl3PtDWYo6y
ypKLwbi4u87NcqTtvr8F+pwIsT6GHNT72giLVtHMtfACbmXtlRog3mgkElaUGcPCSMLKPkzQt5JY
biPtWsCCqtP0RPeCMSQtcjUkZazPxF30adjGFHZVK8nRQ5cDIfcCMJEzSyLDli6lB6qFr6tAvMry
Ri5QrENhm+LicRuqnIFnBwHRpwaHZiXs3g04C+GfTQHj2XDIIP5UWADW3mmbEXL6FjUKv7nWObOY
+bEbI6asaxBRselL1ieU3t8o83EgRsUpgUPY0NGZkRO23rtkvYjAmqYGwF5M/7yvtXOUH5t0plWs
yy6v+sZW8BaCZ1kOfwqimGYT882Cq/kAVS01cCa4P8oK2XCGZt6ThGRs/Ep5P3FF5s4yeycEdo+N
xmiZSEIsRjb3DQWPomtwbxWaFEu+GKyP4CbtU2ZdlUUWjK7ntC8niJIY2KhsnsOzehLAhLVLKRW8
fLMZUerXoZWALbuO3c+1vdE1ZEkIWCbvCCb44PuY5t+xF8klzSu2A7QbMJixZniWazFINlXMGIa7
4fKgDqcyCX/rT3nqDLhoJpL+Lpgp3HMXsyLwPPxsEw6B1VzMoJ1MPlCe39ukWbPE32EULrmZ/rXQ
cFdEVkQWbOvWvyx4x3YhTZMh/q9I+6bIq+jtiZpN3iEQgsxCiH6jB7M6moHz6BOk0kU/uQLmJxaQ
+sr8xCP6iKT8HlebmETHTLGoysdaGy7s9XUsV1ew8vDvAID424ia3HdLZ4f1YU5P+DsbBoUeu3sV
TDcQb2jDMqPyxjND/HEF6Pm6OebFV7SFJd+DPyO3vqR8Ysm5wQW9AAgz/DrgRL0z/+SvuiXXTFf+
bEcGJuReKafu30PngAPBCaZ+s6IprowLSk5KJpluP8KJn/hFNpQaTY+t6YrBW64Ex+6oW+shVXN5
d9m4vQzh5OwvQHlxRjCkQyvF+xFO+3LO+hGi1XS0OTjGxVdQh+BaU26A6jn5vwARYVNV3EDysPrV
uuqBE8S9DR/O06JPasyrNDuat72CzGVda9Qp1ydU/eAOqDWamvgtFROBunlfAE+SzDXVPioScZGX
IIf/2KSkKocWNZ2IYz4PCypvxmmWpbyoPuwTUV7g7m0q38DLnGJucNTGsnWhwkj4EVnkbP6eLuAq
GyGEbVedUpHCK4Q+QkwI3nm+2OInIGwjlcDc1jMhRMkRIksorvlrvDH77s+WjBjLpYUAS+qkFrrU
hElWCaTq63IFzwgUnP4WOAZiaaKEpo6UwjHtZ0avNdT3fcwDCeyfhDXpvqyKae4F9P6Mp5OiKSHP
rhl2xy6mwAjr9dFBZ7I1JlDfgbny7n64T4dp4NL2OCf8Pvl7ElfsaHBYSwiEahypyO2zkP5ypPmt
3zDR+gA0wfUvsEleQxgPQ6eNcXVYQexLKsoPc3rne4nl8EWEQb2jYP8vdZVxOhhTK5d/tTRk34/g
XWESUtUadNncgpAgIrhAjXFXiu5l6WgUQ4tTNzoDBmAE8tJtz/xEx1LKWfdcGioS6ETtObUv+mVe
jzFQm5WF1WPpztEGCxZeRMyHVt4ZqSU2EgV9IajhPwzY/LEeql71taRK6a7PNfh6zSFh5oXQfZne
NX52IxhC2ftBJJpaZ9x8w8TbVDo5IuIIsNGE7KeLVENENxVm6rSEyIpSTkY1kz9W9P1167ipgPw+
8bA6sZjObX9nJYeh9g1degf1pkmHI8a8lrnnVS/yAQa5VO6VCnGC1C6upS/Cz41SD45OMrg4eDqi
bBEGOux6BLnzDBUiwTTUImYIkZia+hrIDaT3M55ulUoa75Ynt9nsdlUHeku4bbeYYEAX0y18yzo8
kzwYJ9i3V0AWQYsWa/K8TI+Q6bLADQLG641/x27pdai6w24K/j2UVN/dqmAlFFkWwIWbx7lM+WX5
DgPG66xPCn1xZ5hSzgojbo+b9QR5gJkYDt3u//KhcN3j8DbEswcwk6CHzFEeJgCqyYgzJS06V18X
TU0p6C2WNbCGLz7sQfrQsKC5oN4eoUODVdLpMatMZDeV+zs8ciLbfCkqCHvQQfXYgN1ZCHE1lbbA
DosO2ccwe0W+R+l0TgSbb2GXoMe27B0+CqhNHyRt1FE7It3vUE7MpfKTizS9YLxlAfZUdhYGaAmj
boomIVfhrOoKTbV+57hIbHT4TOU1Sg1FuvjwUOPYEA3N22mID9kFk5WeKDBGjKq5vuZ5BoPso8rz
Zn1sNRSj6OkvTLzuZiXRXOz6BaRRbn2/kURVjFButfxuxm2hMRNHZPESr9HgCANis19UhdDKN9oK
DgvnO2UjsCVd0rEb/auedRYQTwn1zd8nPtJafAXe9hwsYLS5EABbXEk1wAhVP1+edgOi6exJJrP9
Z3s7UzwJSz6UC6F2AGmcHd1HqbOcYj5i80T5yp+PNsDwkJSu3oNwYJVViHw7MXcEc1Z64TANyByN
7NL1Aeb2bpfT20wvGf99+g6SpBKRGjRVVHo5MOWwk8hg5cgLio9ScbwOMxQ83il6XLiGURHq2hBn
uaLjSTW4zcBR9GkZW75HVjP/xUt1cKEgTsDKBcpBe8GqIHU7HfVWIurTg6eIqqW1d4L1KCO0iNqZ
zo3Uz9S9AvnIw3rZkXS9zMb0f8bdYbHPZR5MKytp7a8LqmySwaHqVxRl7zp3G4/sGHkuYyjRURci
RBF2UiY855v+zyrZimQENDFJHuD86cexgQ9Mw46eIW6aRJFIf8P3kiau7q/sPrmMoJJcvk9fXG4i
GZRE4SgP161NPthoMqNfww4LcNdMpOD1jKVZ72dqHyDT+Eg2a/Z6vyPom70+jcXg5enCQpUEPDGK
POPenzjVFq/N9GIF0E7B6pUmauyWTe8uRxQtAv8zYs1FICppCbZ/yxO7wxPMX3fVnuorgZZBOzZf
71E9qv3FXetdghv/Ak0EGnpvYeXez54X76PqE7R2Q2arX97EKvlV35PvR8kVZZl9p3q2j+As3Ect
RjLubvtv3ngT5Y5X130bDmiNoqCK8MdnTIIbiTJ+vucplruSVvbu0qeTHseJpfi/EszdArnyr0HD
GurC7jQkt+0t/i4s1BiY8QxvdvLOSPXsjgTthkAmoSYK7Cdfjat2kCEolgdmc95cxBBz/OHZ0+r7
OnoclctWvDt6rliOVNoZVI6c1dKdSgIeYOwPwlH1he0a9KXwrmro3Cb+yiPS19MN1KiJPfXMIj7s
JvxUUQSCFv7K6062XdehbGZtBBP7PU63wr8CMd6Vez2eTLDs0CI5r4urDHK63VxJHVA0N9/qidlw
BCu6OtcUZFnMuxOvYnvairZ794h99mMkB1Ybgi3C9yN5G3BT1WHgNUqCU1IL44rY3sa8HylfqOfc
bQWrU/K3hWpLvCG5sgbiwP8ebtI2ofmAKp4HMMdNBd3dgcNETSVA/IiLD0yqxKxj0naqiUvEDarO
y7uiKf82z4+UIFUfT8pg0cdWm2kIi5+wVdrbX8tD5XprdQjuHC7H0BHi9MHSWxJNbaHHM2fZINKy
fP61/dtWXCXs8eLICkng/xqqxc8rmbCQ5E+By6ijclOBxXjgMo98b3e3CNf6T1QeXrhS9oHYG0XL
58ion54ne1qOj3crlBoJE7OjbivVx7jNrTE4LRJP0LlS3rmMMNL17FAQU0k5AnMWfXa3dkjTbIeo
X66iMqO+mJCPe4/cq6ffN5h64tDvobgsqSt6pCiCRD8MbQqU1cIXsLAeqm5bP8Ieetl8zeKqzbzb
TUbQk2+NgbIGafwZpfNIeX85mGQDZtEWb0TVZVtZuzGCUuZbkZdKtTbkVIqu2QhnL/cx407C4LlN
/0WgcHmZqsU3SQdFwIHUtK2rsPA4UGiA5Ks+CfGuWuXUrD3qkYE93mgZvQgLdd7BfXIZQNEnrzbC
u7HpAqh1TIe0fw14KXgq4hjWDkI+AE/UAYKiVYkgiObZanOkaK122G59tpF2DeiHNXg07bBWh5tB
xa18oCAPgGfJJgtb3Y2J1r3SBgtnnfNuFJV0K9WXgKlCaOO7brR2GQ3RNDwTs5tPofQNffHC9YA/
MGbnlUeGuP56tqOkcZzPdXYDzmSAjY/TZDKdkukJli6GQsnN1yOBoYqYt48cw5IsW4qMXrJ5ZhYf
7MMAr2ozs91CN1m1fzCbMQySIcnrjAmf8jxc+sQ8AbBWmKGUxYgisPF96LUtf4jxUZj75At1tQnq
m4KcPf8JS0kg7oHrgKBnsKl8h6uzwu9nWwWul6U1Kvb8Lim5/MMxIt83dT/SjCFqocbLtE5T50a1
fg0U0xFMkd8HgOfw9p7xFNwLQRKKbV9tGjm/fiD7b/s3pGqlFL82GzYFIcf3m6UCO/MeROoGdwlS
klsX/Dnv133Zo200+xT2QZqkVSTld+9mxHPw+dXEr9OMPCIoh/1vSOx2lzIby7wn9w6Y4HUnysxF
vIxqS4rkoftVmDRnbaNHYD73SIBL/70/O91c3WhToonwRDU5HmV9PmQe3PlrO8k/PJBRyOUx0whK
gXP5jWkXrDp94kiaM0TedV1RzKd5CTC2tOljeALStNh8uzgkfDyCpamEaoA8a2HsP2INLDB/P+4I
eKmhjg7H/iQCJ0Z6LEk/qElRH1IoNvPgyL0VJUfBkPK+ygeJgTCii2m/REqPrMOdAW6IdbdBB+rG
qw6gHhS1mwWONuQurpJ1p37zbjp8TxfZJDWkhtEU/f1b2jt+uNYe2KJ4FcflojqJJmzdc4kcbz2H
KNsc+L9yBjOaqM0uTQgkJkH4KX0AQos9UByoruwAVRMnbnb0t/NoCqUm1AtHHn5iwO5DUcnQgiv0
fSldNNOLt+on1O3z1o2We2X+2abTD5UEKPBuzSEIVsqpAcp4OMwNedHcpLBjNPoiUq6i9SLwDzd4
1zFr3j4oD652zEi77Ak8ddzNj/aZiReloghWeJqZd3J0QTqh6fbwaZ2/mjxuiZVsTbh3kFcUybqH
sZNdV5+OZIJRt7Wt92yJmxpEI4kTbW0DLzhPPR+Qu9bQHCjNkQaxaLpNMvA/JNec5//ChHPDF+R9
IFLG7jwzU9k5AJ87qJv/X39xRRlIJGH2FZdKT+uH1Biq05ch4GPQsO3uOpQt/J1XxnKrZTz/2PsT
1RkzSwPKqQqAQXD8UKd7M2YV4t8sTqBQOFnmrHz/ve1fJoaaLlyDWUlFRA1r+QwUfVsQSSeJ2kzi
VdAibteEAiDoRHFmqn0ht9njG1PWxqN747MeLADi5avvxWH+S1VHxxre8MXBPfnBw5CPGUb0cJ/O
nfMZ4WSchCd3njsRTXFq2fHPYJ0XtiJxWTD+0kNKJiozYJPX8wEWdiFCqUfVaPn/fyYhqUsYy7nn
yDToXb+XJ0OKYUyyOsaIz9haAcGv4ynaTerDtp7HBl6DV9DVvP+WY2gayJQdlzos85KiWKxdOyMN
pox2rpsxL0b515yyPLIunWIEN4ORGYb0vxdsUmue2drPP3zMa0Ri3GqU5isoouHkVxmWAFeF1K3z
BHKRxoJzgJfgQ+y4UssxbaN39KgggPnPdv3zwyqr+6Cms2WUoR3a16nNufrzSMKEYEVKojnfgaxm
sj8HfYLK7g2TYz3KK6etAoNGzHejcYroHhJ4mlRMCEjNlYEVwVZwvfmaGy6ZrUzk+PvYzItybLNh
irVFSSf4fKu10dCqaDaaRGyeDBWvWw4Sa1yvx4loCC3KptToKMIKFh2BUuAipHpStau1Kip/lTCv
sxDVrDcLA4pKt7tIsL92YdZuyGclcrJott3mEm/ntbQZeKwLaPoqZNCcOur79fe+Ex/jloEdGZnW
trUsItRyinI0urJ+ZmLQ2kxDlo/VxQXigsbDfKcje1LMDDnPGIhNU+ZSlbz9QA1+KLaAxl2wW1u/
VaLfTDEI1Th7xOnZqPxlIHj+JXKdFn1kFhQb6LFMQq/yOqS0Ivn8MpKMjk5GWOC46T+AFlDZ39Hm
x6OiwbgDtLSIgmWjNME53i0eWPNoBFQvcleNpVPWgZQcA/ldPxwr2SkhIMd8EOutBL5f92H4Q1vL
U1dMHKhQfpm+isMJT6aCRGDwWusMjEwx5jHsM60gPHbFuDq5kZMSfinM0AGA4v+IJX7JriQjYOf2
4eKt2CtggK7lvjoEkjikUkWQdrymvnoAzPC34gqb12wEqNabcjDiqY3fGW6+BpxRwo/dS9l2NMCc
h+kvZskH7MYYRFPpjVIlhoyNYeDkef3XaYFu3LwjsQLjPaxKh6bVxQ86d9bl3tIDCkKyVqYH8MEG
SdnjAS2aIRfUN86w723nTRK0xyiO1ZwDRTFkpGHDR0IaiQxNDePnkl+E51HlNs8djYMyrZDANMLM
Zx26uOwN1RGMvUTFsE7qypQTAA4kowTFSjCIWOBN0SEwLlu0BndEvHYejL49MzsNF+2dwDPP9ojs
LyJj78zHsmxX8xJc6PXIZJdo+guKK+IgJ8dUBSKdKCu3KJwwwXcKWq+lLbtVrV2zT3VVF+GzuJxw
eWzDMAhOe/LPqELgBuUxiNTQWdoh298eS2g6+jqzEfH8pHDbPQyUOof5P9twrBhADB9wvTarlUD1
LAaRJiV8qvqAAmFMqzM29Xpf9md41IXFj/19RKtrQIG2GMr54g0ASUg1/X0a+gqGChkddzBmYwdc
Ev46GAQYjf8iAdxUuPqfkUyhDJtTLeXOblX/otOwY3xPPRs0O6qrrevBEPoA+QHMqTfasX6bVD3z
0/7RjaZj4S0+0F0KsfAbFCWUmdRLTk/rex1hBZZfTvDobp3HU/44IhUt5qDud/+OP7ZnNgDNPsyp
qBhSsLm7hKfBGEU/sUHylF3u3dEH98MYH8xMoo3G8ragi/HQp2IB4bhJBduqoATddiL/KzcFgIk5
zaCfGSb8h0w+8qasx74MeubagieWH0+V3xi3oa+A0FfgYXH6DdEvM9ARV/9qQqL8qqVCNJF4dHMo
0fQyH15TUp9H9MhP/0KDrrPzVlVBzxWGskI2h1vXuyj3nBazZ4TPx3qrsXKOrXV2p/l0a7C8yCuH
kpcPBfO+EuI1F4CcTrVs/wLRmZJE7P4wyCZy3araqFzs/U4/vbUspJOisCKcWUnliSe0lw138hkQ
uj/yqAh83uQepfsPhPe6bfrhVx/QvAa6tyimOmxCcZ+VIVDd8KLHBe6b5oSw2JS72r612Gpoabt/
/5BWwrupgjU2KZiWFXN9wdI8XZL8DYIfst1BZigyXVZ/sz4y2TT4CVdzh5SqhSOyNTVhq20mBRML
l7ga2ibvXUGXJEnnIn3lH2cHBgSrP9bbCEOy2bcRk2yvbmsJMVr8YcaPVkVTYG/efnPe6V0A1rUC
9T553OOc+iRZVY+6eS70x2o+0lFAzSYkO4VZeTOMB3930h9jk7hCGW3IpzXerpBSRmND9kJUHGeE
p8BTPoamXGpJqRiAAGVM9IHjTeK23XsbxhuessYWDd6UhfrilHr1Z+0kqjLMwEDXDPqXtmgPiwDz
8jzfIPFo45pf4/jf8sG/yEW7MzV59eWW5SmwyK5vQIg3VbFe7MbFVYB24XyQhDKZ+PbaYhLlep12
CPIV3xal2f4K6ToXK+5K2/rTte/LaZy2DIG04+ZVaiQKFxAYIwVojDg5dmXGxqbgzeWC1uHnUrqz
30YFxVQYmC76GRP9Cl8EeVxGZg8TtK7EkL4Oc5XA3ryIQQm1zAc/wDceZt+1uBxB1b47pT8i0RpA
9+f2fxlHjP7AsNZVWeRZdiz9qX5vse2ZiKx3LoZk1hN1EpyEPEhLJrRY9RJ3dPXwC0AzURktWWh4
P4oUCZCn+jSNNemUHXV2RbB6OC0mdyf4KDwjdPRdVObcYAN1AeFogwoSJz4+RbKKbvPhJ7tJSKdy
AMs0K+wZJNpNcls9BaYmpFshqbeFVoBupMmgTU1Q8KlMmzsjdEHGic9Q0WaeYGOntjX1vyMCndHI
6v1CaPwpQ6rFKEHBo9zjGYApjtLZ4dokQedmgkoOwwG6+FpY5Xo9OQ23YZjGbCE7zKnCaqEMElxt
mkqwZzM8jVzoJF/rBRJMF3uoR+m7nxQFlu+yJr6uGDwbp7SzXK4AcbeCi7Xj7BOJNRhKLF9g1VMT
dVrozxRp7mr013iQJys5X4patJ7hXcMexi2KKC2gDilMI3NoUx/MK8vD4bBntjamGoztDbEIxhhN
7IpO65FCAaETMls2rozw6nlDQ/0t+QSU3Fv2H1NgP9169hqB8cuPmjCQjbkE+w1AX8aP/RLkLQzw
k0eaBW6gMmDmDx4zg9+PXKoGdt8YbutN8kLuBbqHeJ3tplzVcT2e9ihmZOmb+x07FWsp366q6Lk0
w83Jc2oUDgKuNcp9d0HPpgJfoqKsV8fwJccm4BovgEkjpOsA/NTEqEgnTNqOEwZNHs7Ix7/oERnH
iuwkRkNXv90W5ZHHYcDfW7JZvRwJKTxR9dZjSlKcXiifVI2xEaS8/et9sKaeWjEzTSgYCepKlVMT
nGORX7mvMLVuG9eE1nF3vLQuOeocZQC5GTmjU5sFMcbuiSqVE0BdYNyLyCKN0diQXSjlE61X/QWt
EVDcNSPhC+DXgZ8Qxg6b7eS5BhgpgF2bNt8y2JtFgcitMoWS+pQeJlvLvAlDf9O+LeMJQYkr49BG
h/GTuJ54PQ7lRep5E2WW+7p4VijzNPjSB3fM2FKpVimv68YEnuajpgGfwODjfVuRNHadgC9Uh9WQ
VuO4UivkLCQ5nTjG5awFdX6pds45aAk2zyiM3LBEsq/O3h/TFhGqlO40ATY2KE7AVegHSHY9AnCV
DgCWqPr5yrIXFOETAidIzMNe7P43ZnNTJq7EVHgyTDdh0Ru18Q0zpG1JsMqAOn1ggrEMR9K2AtSv
co7pW04RpCs7iDxGGU3CXeahpe76xXuV4kRwjvtRa1DBpFBhpU9f5BzIarNmB3ES3dSD4ofdCkKK
TJYaz6sO7eNnqo8lDNBRuuLOAgFDrX+OYIAhI02KnQ3hcoEzad2LqCGl2cjkhiI9Q1ZRvnZ4THPP
2KN6KGAxutBuqhHGf0FRNpvrP/sN6OjNzSs0BIFjZBh8z7zYFMfhG0g68uLL6joAS0Xmc3vgVHwz
28eKl/5jmTsNUGHosh+l489941COJflAl6uSV5kNSurCuOH5EFVra1CgwL1AuTzeY+y0cl2GV7eg
IZtyJOtwwuvNP8BYjJU1n023DWw2sY4M9m3nIX+HrppM8jOGeWr2YBMzCMAwBksOyKPcEOhiTNWQ
XE5v5wTOS3xWgWgKsX4jdK5X++hEGao3g/za2I5yNZ+9hciouQ11F5y5q1XXLlHfNaAaxvfdq9Fr
dqDjTuN7m+kSZBvq3akL+sueAS0QClbrHarcIPBUMPY5+nQUZ444t6e8tJfyTNxRQkLnFkqAq1Ji
7XZghMqXANicKnbcSwcnXl/qwQ6hAiWsy4uk+xeJZZTryS9R80E9dewEdFZPuHhfNWGhlbRiZvcE
fvc1IKF1Chx6WMWt54Ok+zmVjCfQkUl6Q+8vmGeeav0CqyyJFR4bEH8f0kbDNuRGsWOyf5V68OP+
rTmw1x3V0INkUjaJftJwQNzkBWt8C6iS/u2Wd+aQ89djGjpG7h9ygrz2d3CPfVL8Rb+D06MGY0JJ
B7TLa6mC7vx4vWkZrmwkF9VGQTr1xagWRbKQY10YyKcnDyVdDClahou5VyItWOAirW5+sZY/8AWD
UbcoEQDSInK8h0ecnB8b/n/J5iav2V4YWgt6PMHdnQnJXIn5eL7pZ9l2BmfKvV1ew4UM+6LDqK3s
pOvptTI2J8nVTnd7XAwfVj+Kq9wen88IJwTO3fhr7yffduAQ0piNQnEXeIHpBeKN9TH3tYcE5zEC
tKTg2M21jexFx5qAMHsU9O+tVSgSQXT68U6Ef5fQlSGR2/kBEg8bP2Lx80zRW3vnTsq74i5A2Qsl
CwZVJ9/276Yd5k0RmUthjkrF2x5CPnvBqdOUCJ1fyH61SH2kXAG4+b87VtupX+62mg8hK9xduKQX
z/spQ8dYehf3gswDBl7K9qGN6QJP9+0imQ49nu8msQp12efRAWRPwNY/m3cu86RTKvUw9TM9G+vm
++aSE5dKEbLl45WiqLo/HY/LFKjx70s5OYg1A4tV+aeApkYsHS3XZ/yKxkIZqycelClQK9HuacOU
2EMhoXGbHJvGEUjOGyB/InN5FLB3Q/sy/p6+31ZUm6+WDD4Obwh2SeQu+XZLcCdY40sHRZD1+FOe
Oq70LKagHvsK9Z+HLdP6a05dz4O+aZkF1p+45432tMbk8T9srWQ6Vb65oG3FZWXsNm7zghS1lO28
Qz+4kaAx3VgmBTKl88PUbxGUVRIWAb5DEPizWUFr9pKUq3akrPDhJBQg2BWcfdmRzsA1KYfKtJAh
N4hTQ4TiF1Wc0ceGYhlDCwC7OtFCH+7yKLh9/nqXoXcumCJOG6KxQdNwgrcPjXLySt+oliiVyOoz
kAam0crlScyVB7dQyM27jQyq0/aGkNkVv5EPH5FpohJ9fOXn0NmxdVZTUl4c588Xe9DYNFjzlR+h
Edli6M8LfGZzeOZG+JwinjjaPfVyMWRUeAYjU9Rs5eaE2zaV3bBRm9323Ti078hylm2IP81wlDmX
cqTDUscTOSaMs8qqgs3l3bG/0LPTGtqhustlPLuduqdpPvAws+Os+yx5F8paw5NYo32oPlUuk+dN
gVeM4L7ZattUNjHdp09uPF4XYUO7BgWiXXLGjVMUSLClm214Co/jgA5v+w+IU988gOH8UoZMZC61
jNC+is+YTebqxc2eSUhaSvjrE4GXSw3F7Ps4Ic3Ci0YEx/RowcgXdJFs7TI7M01z2ZdCFV3mXLn3
ABcQ6FNiSRON9j9NXT8Qk4jCjqzAr60vbZ6L5zCQQSzpT51AO0WlPRHz1ktz56T4yogndTsgYWZ0
eKkGYsHzJN0TBb12YRfsKfHcG5RZncQIHzY00x8mu6Ut9hjo+VUtNnHjdt5oVDFRDVhZAuPQ8dx6
W4GTNvvD6wcd4zhogkeYDlA/Sqm2hw7Wj0v89SwN9vDfw8OWWYg7yPaZYgoEUCeuIVAwZFW5QUMx
sgrVIWYQZwvPZ1OgZnF8H/LIY0swYyl/CkpRZwBSCX6yx5avDOFOphuEcVGXLMa27a9slTSLVW71
MIKM8SdvEUYtLyMTCnJ8c8X3Pf8xh3dETYl6kXGO/nRpODlg4n2JsX/rWAGa4cw+vjqwu+2nID5J
EGsLB6eM6++FENLMwmDecIfEOrEAMwIDC9R3fN0rYb8wSyB/yXX22Pw1RPZyN8+1vadf4+OtF/Q4
Snr0zjMULRJA/AImFGjTcthwwT+/w55DX01aa3KS5fIHoTF0GjcWeqxtJ0pTVW57UwmggeTP1mVA
1b8c8zggj60pqmwK61Jym3l42w3hD73lbaTXJrK5Wrxuuk2TjjhSDS/dXNpNliPncL1g51C2kVwE
dqTvQQzFrR4T4S5XulQOPAEQK/2uxhPPBAl8zVfXYpPuwOxHPDNA56Hw2LqgCvDJh0/hzGysJlts
ptFnu2AvXJRArbTfe8ZhTAHaNsqs1llhxUQnfOXz7trRmJFtUbbskFC4MNNZA79LDj3/JIHkG9xB
iQ2MLNkZkEZmkXQ/RnBNNfJY/l0jGMkfI3wCwp1IKE5NIWE4a25v/c8pKIeXPtTnZlLlcj1hQoQD
rAJ9Ik5ivfYEKlROeAzEocxqpK3wVUHFcjOkGHV/ImVXDRxiGKoeEenPVYK511qyGIUwGDw3j7ih
t9kCBrXwX7v9vMy6rOK8zUbnnId4BwnJWAehaBIXfGmKf7lvjhP7V9JaLu7WD3yTELIu8jdTJaLG
7PcS700RyiXTZQXvJ7y2oihX7eJU6/WS0Yi+pgEwFytaz2sw0fzUQ7NkHTYHsFX7sXJ+iXfe74Lw
2iyZEDwxpKic6O8Urss5KHCEHGjXXU9hpr888oxDneDN4g4wzK48DZFIKS5kxlGhNO96a1oQc8R6
FWmRFfHDT2rLhH5xwv1ZEUlfK9B8Q+SPGAONHKYRpnAGTNr2qJj5gRmVP5cxZbBFZ8eqf5aFIQWV
gDdxo8LYXKihC9M0Zhg/d1bvMQXQue8+uQ7YC/5TwpnxkaPJvy0WnsUYSBlTzkw3kMCvo6a89oeu
6R9fSDGxfWXxqS7HsJAeFsN6ZArsEhzPp3i5yfOgIwJdRNtiX+AOHh5cRyYwFDSmVKp/eSlc/UUO
bdhp/b4/bUMp0uvKr41H0pyi3pdOGZNuP78X/72t4fdQmDxomtnZHOszENxG5J53JQGkUknxuPG2
2rWVULH3S5B0MX9fTP5odB9p/I7oMmAduSiKhO79uky7xeB9bk7lMyiBjQ+KIXmR4kA+2S6CsgZn
fTCYyixXQTod0CyEgA2j/H/WosBgIdnEIGghk8ipEvXW7w3ecYnqzYNWeQaMF8GQlUHx7l63x9qd
y1Xagbv+MFIrW2D1MrVXCTpsgctH7tS3aPcfwTg+4NxLmzuonbPI2ur+t5KiwZhomVhvZxy7756w
bQ9K1mn3W/ZmWAM6Yn1DoTa2CbSWd2YEBHGB2O8DsVbM9P0kuXOmnIULEdwRDUsjQ9YzIJYE9fut
tGpgjNzMYZYiUZalDqIduzhRfWmmmPuQSLUzfbBu4mZo+nQzRgJkNYQoT9woraXUUYQUZoMKMA5U
L96g8dAfCZ8zyZJmc8eWf9YuEa4xwiKWZ+7QZNutWQMq/Vvtu4Q37GkHlrlyWhcYR6tdMlLYWxZC
6XM3pCApkqFc5vTtjhgj85xUEKX7WbWJLjXrtsURmDbI+ipWAxiP86ZBuJ1NpCYBua3bHcsijaMR
uqD9vWKlGbkI5vm5a33JBymOl7FzPD0Oi0ZHDMpBH9LJMeueWIRuXvLHvRdZiN16Z9AlOvpLm2z5
Mdrn0ACY3QHqNtPo/Wo7gdgHGU93euAlWcQKVbYiWjWhSUqGEZdne2h3q/Ls38+gAK1XK+5fPCOz
24rl77wBtlGBJh/CwE07eYyPdHkGQ5G1tPa3sK6xvANK4AFKd/1J/KX9eZF9zkMI27+8girGXJvc
OTDd6PHM9AU0Z+3FbU60B0MidmWOjItR9plQm8a23Dhn09PiqeLeNDhRAndZNTW5RnZcEJv7b3Ob
f6JhJ2ZgpvrQpBHGSwBrT183Q1vUIgeZB5lTxWhaJjIj+gwvugpfNiWSC4SjxpwTeA5X0KJeFx9y
JFvtmW2JYvSCNQZMkgwAp+lMMhlFs93WpHwGPdC3efcwxkQRpvqckzY88U9xXv3SRYzX/+kL1wDg
YWrgcSOOc2+4kqzSv3HMaOFQr//s0+77bNYGb1OlgHIzpmk5IyBFpZMmlztsI8+re7hBpD0MAr0J
+hFQ48if4zqi0dm27Lvi76eAlvP/kh32hR3fMr/y8AxramxvTKebemo2TJY/e5kS2JfV5FaCvteH
9SEY3weIAAk18CfRp+ziZGgeyFkf9HFhBs9ZSZ21QGzsfJ7edH7E5PU0eILTIAlwnbUQpBZwnooK
3bNP5tzrnssKYjmmR5XGvvbTy4OWSEd7ig6ysw+9tRQ39LIgrlAdDX7UCNRG8Ppp6wJcaAKjpWKC
uL+JtpvNn0OYf/28KoB9/ZD++j3JMzYbMiiODcIOMtE98MRdJIHW1Sb/B6TlnV/sfsTbYtNS75mx
ZOa6u+RUsuaXIeT9+/VQZZEWeJ+Ffs5vANEK5gv/DIF5qeocDzTn+DxwuyTS6Tc5SDWEzh0HLyPm
hyDDqajl0mEfk0etuyxT55FFUA2tjBJp4HgEewMKKd0IAocKR92ej8vP29hAlvItt5K22zS3F1tf
xceI674jKCQbuJ32A+WoCS2Ml3M5qV7tg5lwutYFGVIhUesKF7vIFpxbIZFxhQti/OHRGI1S7bLt
aTB6BgMPMAOKKOsvhJjALThb7ilEouYypEWtEjLdVVPPGf5DE4vE6mWLvz4U8gSm5T8X+im4TFtd
x9LqbwE1fPqGYMw9V6FWBONg9oXPPI3BvLHJvf24OOsAmFNkJNGcM6Z9YtJ+a+OZR96kOhiL8N2O
yMuWdB5lZtmEGC18ztQjgO/NosBKi3kQc8Ae2bbyN4g2+F1r5eh7F5LH2jZPz6ZG31A3pEt9PIlq
zKO4zUAmFoT10ihO9QoZg09wjfFCRNUbhukzRi74mDVtQWLPqSUn8n9Y37oSmEUJatrNY8kIS2Tx
PVPZ8T1/e8wyhGwFlOalKZLJQjYce9i6k9QA+k/awoUviflYyZbcwT4MQhZqVbL7ew5MEcAdUQQb
MOF8lcidmhheLIfP/Uh60zfLOfO3c8dGKO65B3BkTLq8nz+S1k1stQPa1mQNLqpZ7lMoje+5VBBl
KiTVHitlKQEJrRp5SIOdYlTHG8mxdLL0F3Z6QyIFKOmJ2aK2E8IpWyvtVznWt4q1iudt8RICPouB
4nX+VTtxZgacJBldHYStuCLjusfySCFi1mfv1phLcOOmufZE8DTbl1/de/+/6NT5ee6LYnB1K0zC
WlMyoGuiihe7HajRbMRDd5KwfjV9M897xKMkRpU4eZd8xWg1P6vGmpTY32iQ52Abm27Y6EP+KPku
dsgV82uENZ/J+O4TcqUn3y2X+TQKLYYxKnw1o6nmM0aLIbEde/XisX/7sUSUs2UPbcdqqffbQXbo
HK8yBLteZtZpoYyNE2L3QN2NboQhF2IwJ9yIKeTa6NXHhG69vOFZjNjCz6x6lZEklisxwWq4Tda1
qJn+36ttGXrsM3tooypaHlmGMJ3lhA4M5ltoi+JGNHpGOiUqK7cv3vqDTqBnKLrvuN2aVfnpeLSy
RPLRjICkG8mRNSEoeXYyLZRMBjZTyDfNJkA5HkYgW+4aRMXYhpzCwH6ku9A0Mli5eMMICn+zICAn
Qi85EdMrQ+ZDazSTCLEv6nJsVmAHDrYTbNMquBamFiC4ygAE4Bph3rQzLB7PvPOwUjNckc369LUx
3u4Q8diXFExcnsC5sx0z1owPeyOjLugabkSRQkLA2KawDV5/0ljo8E/yymDSxY1n+U5ysk1taMaB
UCXs03mUEc6qNARLvno9MVngr3MNw0Sav/MmwfmK3qubhI9aMAcprvVAeG5SDk+6oB9zvoo8sAFz
7x+MmE55VsDb9atUwGdGyVjn+zMQUg7mgRV2yzIwVSk40/N0QnP/Y5vBWSByzC37ZKuy+Uj7KhxX
KsSc0KxE8RO2O+Q7s0lexLhsCSp66HaMJUiC2ZRGCoPvo4VAyOQqzUWiQCplmm5tJ3Hbf4Zqe3Bu
DuCw+dU320ZgYTR9+xdYDP+UKqifft2P7m0of1vjPnNVB/yJiXrYbZO41FBPw1KfyC5AQIqXXX+M
McfnWTpjB97+lZVdstjurI9n9OZ1Noye5YYgXB9zewYa+WsGFDE1Uav1U1nVkBagNCfNBcsifeVy
bELrSqP6jv5Xrp7nLTyTX5UxFj9XE8ULdMooK/Eh6Zd6dTrq4m0MdEpXZOde4l/58lCLXcNfJNzE
lb7ta7nCrr7guaOt9WmBo4DOMeFsqp+UojiEqf5UDeZAGJpcmUSQMVytkkfGnTb4HGcqPVDNo07q
667sz/5X8NzE6eii9GK0xaRr168gmqdBqhhgmf6DZ1zi2ZvzUUWr07wq+cOGqVhXZtp/GbtKklRK
9DPAlLaw63cGaQv8Yh0WtwILGB1C2r1NWeYxvVZQLjwfRltK7a8Q5CWNzNU8heiDHuGcoLMoJ3dn
s9nod2CuVL3H66tBVA62oiLpT6cdODB3XfnH+5rdcxNOfGgk7JPWRUcwZIqB/3eIvb37Io50LsWM
EhIArW788WJ4UyrwsYLQOaN+0wrKjsFdsxD09wAEMK3aX+orUDwrAz6ynTgKy/G6bTkQTk2Iidzk
ZpBBpcn0KSvUd+P16Rg7KkrD7mrixFLJcG3flry09fB/7zZZUZWd3EqVG5qU1XIs/b3rIKZggirO
uxVwhzj4tqZk+R7iJZBnW3IReT7TxIRhKpeh1W2HxU6zDo6XBF1P8uzoPL9V2KdTbPgBI4LL/J8P
0zvXPqQDdDkDANZ0Leo01WwnqI+g1ehG18uNgFh0wufeenQi4g9H/BtZvic9wG23Vro+Pz4UCO4L
ZTYFGwCdJt5S74j4RD9AhVnAdTF1B05R+Tdxs8L+gWMvmCBPOamLvCKnNF1jt4790q2rFgUMIWZa
Y3mkMDBW5Q+Gl4ItPrsZ9aWT+96v2HSQ8x6+U+M+kmxLeHULwEue+ufedh79hUbyIg9o5iXii40L
IZhODtzzUd1TCkgothitR82m3QH08gt8Pd+aWTMCqOSfe8s3anWtO4PN17TBENgjP1VzA1+yB5Dx
/MBR6KhkPphfhlW43Clc/9n2kOy5hSglyhHb9GpZEY7Mbe/l1JsBIOtrWwnOsKXNipMnmwB1EmfU
RY2z9vsYVEb0JXOg9xscj05+pSuJ9X3IsLErqVlgmQb5mLO0kRxMDMJaN6+ZUBxem0tyDK23n3NL
roj+oCoq2YbutifURaLyLg7xvl+sOzmDMpnVnsabKwIDB/MeDWtb0mrOkhvZ4HZ5ErNzDrRsP5WK
dczfY8dj75Wm55WELHky+WsNUXe0NVsFXG4rzx7FTr0EURsvJOrb2jt/7TDWX6kZsCHscvQMfwQk
gXzkOpO5ukQkdmocuSow3Yt/nLuLGKOcYK5riRfcmeRRoE4a7u5XWK7f1ztZ3y+YGH4DfIAMTzNS
QSC9F984eNpSeMc2lNCJut7QyDu3nVnnEg2Ccv9v0XyqsiRipuS7xNTXv5NekLZHcpQZuHXierXx
rDzb8YBa7aNVKj7GAPyg+mQ5GwhQmQzYAxDG41+1cPRGCxPSR+kONg7u43qrgGxS/dD5h5lQ10dw
7NqIdIPfYkfWMDxEAowCCT9LjQTjVRTJwH3O4hbg2H8cFTKwkq6F1X7zSROrHvdONTSzjV1noAod
OcuA1jMK6ASa9opQ20uE4+R/eeBEsC7SrGB/L48+dg9pjlx/ghHN5hmkyPM9LOBiXYyM69OJced+
ywVzAP/SRwk3umGohfBtjtu2PqoonDXYf1ER0qhBhvuOX7bAj7fgi8CQe8VACewoAUSiB314M1N4
+ArojMdLVvXr8o2OiyxkJD8ON0nT+mjJ6GSe4Mqc2CRW0wWO7ESjFpNljFe2MB6aXDLILyIP87rU
BcBAOhLZtlw0cD9U60ix3P9g8YbxrDtvmrrQ2kikcAiBdCXlQegp0gjh6mI7CIIx3shvCcpDzaXU
3YVVKV4BLM+39QtUeFUdpIUeKlt3I3suuKptq1+cduNMVTj8V5j+r6tnpDBILe6F5/t2WqUYXyHc
76hISPUOCYQh7wWDr1nZGrZ9+6jAs+h9lS14ytqCBxO4DJKS5R8oFM2Y9vGhLge9yp9LVnmzSYps
l6be9CkDAvJaTsvQucrdh7je85TvNJ1FM5cOlqcdHGCi2bUm+N5ATKoUmRduxY6K/hqBxp+pHRUf
kE9DnB7KxmZuXu1KpAotrcjVqETfX5rrUxtKNNEZqkWgV5Re6BsWb0dhI9g8jJV07KQ3O5y/2+J+
Wlmi1dKDNY0a4xq5mSnZxGgqCZOu2pPcF4Lp4awUCOlJVOwv7RgQ6wROeRp14d5wVXSdaj78/SI7
J6UdCBYtt9n4ox5qI2hbG2YPE+XvFcwKdws5+vqXt8hge3EtIWsC1cHJ9WtZx78Tr+MPXqi6JsHt
t7H5CsN21ftqfjGZabG2fW3ZsUoFmTgehNIBTx6xOYmLLWovQoQ6fJTi2GPKA4FH8c9P/84i30Pz
cB+2gEC0fSJX63f+omW0cBrpZaqxB9maomUwem2WnBmn+uJjAskR5BaIV0w+M1RL2snZtg+y0s0k
RRDXs7nRvV0ZJvtSvuiWLutjhNi5RrxY0h/9cPwleWkQVfRNojPsruFTp6Zas9BYSrqM01NoAE4L
E/dC6HGZHc6SPAzpXyj3NBSuKDcBadN+r7MHQLsK6fkydmJzVi0PukUKW3nR9AwaV7ZW6k1gZRKq
LV8y+wNXoIPlhTPAcaBnKFb+zQESDaJFIODMC57chDz/nWxMqRew9xyQCZNTrdB8/lFgYb+yh9FG
V6gHXFiNZ3E1VtsodzaOyV9tZ6HU8kXIkg3Ga508LG09nrdInIhGC7ivKHlHqIJtPOh8Hb8JQRUC
h6DRgOyDqXnj5fqOagLBfjf0DN+N3hZvtDf6Z2DGAsPdbA97UjJxAT6pQwpv+bqNYqq9uiPqUB7C
UBFz9YW5O/a6hHscJ2rfFCsDk7Nxb3fak9gPtmfHIu1ljwXjfoVh9DN5i+zlprbRlrYHibbW19XG
/POHeVBKvpRu4t5UQ04QMm8iB1QSP29Hh63exC9NoW9lf5Jp74s4Y/6FDsKcaH8fse6iePTcsNSI
7p8nu2EwTHx3COPqumv8Aspptptpi830FnLZWRAXnSt7jBsu0+Ww1vHlHGOwERf41qDhF6qkc8+h
/KKu7UZeHhH9U9TsfgWUuU4EXukVDYgNzwEWNRTV5gk03tto/YJ4lg62Ng/8jjj7LfrMEtmGu57o
s5KUYtnNdT9RfiJidcLiPqkBWzBrtvEWw45/R5/lv7vDMVrQnUEn7kI8g1IyaBadLwKrBjYorbq5
CdNU3HPhdeZuKrThzpVij993mbGnrfCW4iDlAaqgy3/Be+vVSaa9EVH4yjaDZ92MAl1o1C39JmgM
r+YIyIw3GfBxjK6PSiTzFbPDcpECuLQfgeBvMnAT+/WKQCcFMbNGQh7N9VHgRhcJTw0re8aluTld
xEkd2yAE3hXjoQgsBN/b6zvkfeb6vVBBDzeb9n51IR9iB/DgRzig6xAzYyaGU+oFj32XsbVCuHZh
kAgBeDQLAz8PoOev0mVQR9Ge+8ez9mUmfbLsw4PJx+rxkwkz4dccFYtOGxYzhCACR1t6ZS72dXEI
l1J3uEbhrpnWRKH+2GX9nrp9UPm/ity8Q1jxSKGPgIoh82tCV+4svG0E2UKmSHdHNVThOaEMGy2l
6Us5kjE94IIrocs2pj57A4ZwW1UNJzbGO3NHE7n6mm0p9zvpTJBQ+usUg+ONeASIVa5Fljl4T1k7
lGP06DqpGodcuRiy0Wg7XqZvNL45oMKRVM9UM8JL5+DpD7020hw++Ln4Pub3s1Hv3FRfQ54z6MM3
nwof/6a6294pFGh99U3zx3B9WQRdxMHOfA1i5vvp8OtUUxVlodhNthGpHG43etlc6rbbrN7Wjdiw
6KnSv9cOiq5wACwNgOQLtljMmRXCT9Kib0KolS5yL/FmskCCYbRR2oSxXGAyzTVxU6ZOpkrc7WQt
SI3e/84oLMWHQcITo7Qq1yoGJDZhiwg23ZtFD2/0nl+fYYVXRKvgqEpjJjboUsXDsacA1OKXZlp/
LCEsv/0hPZpifEwCXrpD7DPlz6XvkPRY88GX8QB2c08gMs9sATUTCNRwBVA36hvl4Nbl33EpBoYA
XJ/vbEShwB6dMpYH/1bM20D7/PM4OW5H50z0P/O6S1oxTnYJqrObARtrCcgdodXUFqzchtIsV9hQ
aZHeZfW13awsoJBVXT4t2R7nIUZlkbFzmSpDcUR8n+hRTvcnzqLSdVwqDGXcGSJ+qjSyCTu1A1xx
nWbJGFIVRQhNHfL/XJF8wFy3UJwIE8veK38F0hQdKyHQ966XTT58IM/Bdeu7XQhDZ1eWpnUTJXiA
goazpyYDJQjWX/j3x6s7MwKLGM0AvhELIpeADsQ8n0B3Kob3hocH2FM2OjQOJkm1HMxgIVxLqD8v
RCAp/xNHXkOXeBh6qputYy5eNiDHlVRl14Pg/oibHI6MUx+3koYlRbFJ/khbPksTcWxpISHcI78x
mVUwXpgdttNaRSSxXhsrTUM5Xy1T+6WpRXnumERKby0iP0XVCT6hBgHVoP1pbLPEPzU56y23bcRK
MDG2MbT6aJ31holPKx5VgRBwcmucZiUlspzIOgjODtYkuWaU7G+2BCezUE/y1ywOQHw17D2FliMu
LEQ8ODr3SaF8691yy/synB+lnigl6LTVFrUOJKg2jW+WG7aUDrY18TdMzyFKolDL3xrsxRDA1h7I
to9HDbZRz/7X0lYEdAHyAWko4tWzCZyX7OChj+PeLBrSKzKsMqKsaYyI/W4MB6+UPZATp14Y9jYX
PANWbw7gnTx3H+a2x8tX9U+N1ODzYkw8k5/pFmI6ccmMDMBXJD/2Gj0BKzq/1JYBP+RKr9ZcLNO8
mpYrjTEVsDW/GaFuVtFxFnODEuyOCMwbfP/LlvnIpFgpTzk6Jce9Gc/sb337Hj7uOdmKWuvJjYs4
ryg/2UxLACWvpzc+6VKuDlFlMiclNG/M2FGDGn6E2cz59586p/1U/WVcr4YZlAx5PmXzC5VDoUip
hBF3cSSPtzB6nL7RE+zXHW/T8qI6jU5SdV8iflKueNeylS+lw7V379mrdb3USB/FRCV3GWBT9FXU
NhFSNuN/ceDw0DV8aGMGJVXwManRSI+PJpNWYhuMAHzXovHhqEr6apSTgI0LNeU7ybeBTmHNsxAq
VmUd5JTpb+B8ErcUQ5uvNB8RjFCM7r4czSuxY7V99hQxZdqH3sJRJTA7tKKq6AoJpQ+DtxIffJWN
rnel6TQYFKxmI19oFQ+41wLaSWnaEdkn1ZfB+IhQksAAGKM3UBe0NmNROnPelZV86Z/UHo+jDsu2
nUHiNSBhC7ktTg2PXDdw6rGhO69QWn7mdCAFWCBLnvo3plpzqVPOxJINIVh19olXmDcLrruWUqfU
cYqXb6vQSNWMYU7NISVO11jFqtE5bzypb+UvmSikGJM+cYrwnZT8hZW1UQ+0Wd4/F3OMejH56H+2
HKQ5e+HJ8zn/UY3K/d3DFlwCzUaZKXhGgzI6SoO75j2rxcAOtiBkntbCJ+9yCU1AS9K2xmj2k4SX
lz1c+UMZ8Ouv1/aI6jJSM5O+698BlQd8kHvpmaAYP34l3az9N3QBZ76GMsUrbvqhk3OSpcCMBI8C
Xlr+XoPA2/fnq03pObWe0DNzwXEv/YQNO/HFq15u57+3Vzh0cu3lmho3V618nuL6ktps8zG2oeUQ
v59scerkHBrYTojmWGLkCO/af0/BOhIjTfWjrHNHm+j6FQfJ/isi5f0gjlNSQmfnjvfvBCxW9gV1
6f3dc5NXKNs/zTcrijJaxi65upUXDE7EfqQ9d5KoplnQPxJGjuEKVyke75sLbtJZjz2SsWE5y9q2
19KdV5UvObsDT9ld9dnpwbMevEiUfYbzuAfagbNxT9m/6HaTD3GOYCVDoCDv84/231itz7F3rCpu
h5oas5tCYW2dKhtTw64xn/+4PkAmvSPZEB39QJr3JiK7D2m3x2xu/CQ+lQqod4LNGSLJBrFjfPYw
tBlo6UeGIMDHv9zmpLkvXVbA+Lp8pPxzPQVAVl+6ykC5NS5HZWViGxdI/hLerP9sFbo5f6ikpbr4
Bjy8mz38n93aH4tbKH2IuY1XZBwLJ1urgjdOBXQUDyiBZWu3lhJGSjSrisD4XKSjHhuTke1LQZS1
80E4K2gAcFS9+VRk3IYxXVxYBKhezFe9Cg+uPCkz264kD32f2+8UoKtsNBEEdPKxWKPxFKv5QAIs
GGSxEriwwjfA6gDK83PzdiQZ3P4gAmMUsRlu7jL5o3wZUXe3bNOjeEGc2PprsGTWWI5OkxbT8juF
01OUmEs7zwvs/YZUfdFFhk51C5n+++atL8/pk+fXrIX3zToo815S6pr0NSo6iL2ZQyB99/7pcq4A
tSV/Xi2bbQf8lQWbx28/DCE9LHlNiSm/56edL4cPbjux5PQE/T/2CRXwVIrkvw5d3B9sTK7ar+lh
W4Yj8JOzFkYSI9H/CegKhqvY7nkc5ZwAXxRhYhN303v8aEbBP2vAT4OxO5mtVZXOPcBwOimEwAxg
DZN+WEJTZs26FVIkMa17LIYYkXlr7S7eYzgtCwvnJiOkU0IRFUCF3//LHg3MJM8sUOsRDYdsjs1G
/YWCjgyfuaKzoaWm/zBOZJylOaMmXXl4B1gfBgzR9YRQe/TpLCqAS2YVaN4YZt9LXrQY2793wrpR
T8nn4FuF8O1b2hlLfsOxlZJLeYwcugp4o9PihfrKEA+FjON3TV9RMgl/PI2C7Bg6W3PGJndR1FdH
nkwOgzbpPSnDEn6ndpjRU8OmxhRxU/ShiZf4AjSdyBlJa7xObtdSmB1ae7PddZCdbisoiDdKb5OF
bKB+ssBKCRActUzUl3aaeTHi8L3JqLzcExpG0rzS60PmUHrVEUWDMXFPHPI7/fTj056GLlddrMhf
tcLW17JM2gmmlN2r/VkT3OHveAMmdDXcFpdpeiQR7bXCtFO6C6ULstl+4zmdEJzOQTJtlSgcxQVX
BMEGmGhXjyxF/hsc//bITFtSnv0ZgG04E+bfjmyf6pElfT/D8MoS2nPvxOezydGuuG2AOi+JDJ3P
QR/2oOugjZHq43wVkzI+L/H0twBbqWJ+xu7sf5g/FyfY0KAZDoUDoEudgVRIn519G5kZg+xsT6hf
ZhRUAqsfisySR1y43Oe378cLKWle/7oIfE0INWgpN+MP3VxtHXWKqJHurG8p/yKJAI1lUIRYNgk/
t+qq3AoV6ep08qrXHw7wMPUTLu+5P+O45hbnGGbeFVM/vrBT7hh9fHlpRwBBVff6G/gXxwgnUwAI
LxJA3XHtEQobaHDHWqI+7TsUZDuIwv58/hz91liqX+pD8sOcX5O9GLkRXZoddGaLlgefYu8MICNS
ihiLoBClPhfpaoEQfjgZZchqjqTXyRmofYfaP1Sh2BoApz8Mrg2L6qLEFDyDxBeKPE9NaXIhgz7D
AeiDIXGFvT4gsiEdcrGcP+UNxbVsw348VdweFxxfSofjc5Qz7ueWCcOnI8TUxMsZUmFio9NLJTl3
w3iMUCA2ErJlkCx39m7pxSd4iCYD9vkf1Y34kY4GmfeoLP2PTBELln8ZKoFPfV23F0gF1b2ztKxP
nHoPF7NiEVzswbxUHc7k5uZoCD4f14/F3SirS5hWLyBCx1Z+xHdujLI9brMkqm2OBMwnPqfTJXtS
yupUduPKgDsJRQ3qBTO5HsgDbU2Hy23NnZUtcst49D5S/SCGNP41Wd0KkGV55j2+rqZtP8fdYbob
armbBXdAxsUY+16hL+fpe1t4getTvbHc7OEU6th7F6XRge0qtGBnij8pPINmKoeRLEUir+RvoT5G
2+rbpCmzsqbLX+1gICqmO70u8WnxKFgsqTneYoBcnHF1pHw0MzhuTSMnJYKoyLVnfs+Ix3fpHyLv
jPimUQTTuL8Tg8hjD60fN4hcMFfGHW0JJI9FI0c7bqYb3gxATgJvMPex6/M2+/ecwHMcnpT5ypXD
feYvZEB3X9bSpSDZSvdwkzOj+SiDmPO3AeV3GC+SI0GWC19xV9XKRYujxdvQRp0sB0eGdgTF0F8I
97nU/1eCLS9LjlDlGk83vUzXHbm8nU67vuRCwYC2F3P9V4iRz5I+lNtdwiGfrz2ZO0Vq2OdZFbiw
X9o36DSSvFNPnZAeo/Xn8jEDx8T4BzNxhSzqerMeZDvzdLz7CpmkDbiG8Vof/3ZsUHRvYt7S6aoe
jjyJ+zXuoO/6wufmWbnGemtFk23+S/hNOaHD+YDV6HebqhwlHup259+zfGb7cHOrFBlU5xz6eITt
Qtl05bnpoSMNi7o7BtW860xP28Mwg+pZgB/YWGpVKuL2PIi3KosIdjRDmQrBPdtCpNp3XCwtZjl3
q1mHAbHNUQWpmQlLrgrPNFXvDXQsJHl1Q38mjFkwlNWdFWt9YG6GRY/TpVCnE3InQIYJWznJM7yP
v+8TA6Oy/SD7MUr/C5OGus1BkTYqlbkQ91qlKKN9Ha1ocYLiIZSR3mHkY9fvllPomMeWdRQk/9Fj
h+P9HEQYd3D0OOsd7C7GBznpRMETV/rHpLYTGDKe8XnmhsQYxgojls3faR2dWIaw25gqULTafxp2
tSPq7Tday3do7RKaOMWhhHy9raed6azNdtqWDVBKcxN8L0gwQ+o41IT2BaG2pJk+x6fzYAF7Vimw
gM6Dljdtu66Gvt4614FqMWB1It+wo/bNHkSCNtIKZZ7a7NCKGbMMwm6MmgvLx2+c0glMuIvrohWc
pPPmMjFn2yob03EXdjg9YyFgnLJDjqoXMVnfj4jCquFxRGpwMBPjya172inzDOtpyWK6fZS6NQMq
qt49S4CB7qKh2R99PTrCcQHWEaZ1f8IpKYUcrml9XDha+3U+SyE0pZAlg8fXnOixGap6gjWIZSiw
VJwglDlZd6k2Fpt4FPoRrWCV2rzhHi9WDD8lTNLG7pdvWn1k2D0axGsLqkznDJqZagKeYxAv3zo2
sbSxHIpfaYydrmuc8eGHIXfc4ufs3sQ1m523CFcETvtk/28CnGQCBoKfwxJI/XYqnazXyDl9icn5
52nI//g5627x+PTP5sDaxa7yyS73/r4gRa2rUdKxDBNrJ5bA2vVJ9CwJFbox/N1koR0ucNM8HqyB
VF4zWkv1dj7Yg2I084ZHwVsiORipoZ2O35xPI852Hr2dJHlMD/ZD47metx9ENarFYFqLcgUY2bTn
82oYAO5UOz/KwAE0On6UlTUqFP7D72/x/OuoyYMd1V904+7O9Upy7AgvNpIXTs2sqjL79/D/60lL
jKyX8oHBCXKIi9DFKsrmB9OGnZkrfBH5CHFW3ahElUpi5exFsYiEGNTHlBQh8ciyTf5sPaseRYbr
KBdlctflF6hFrXNzI71SzlBzHs6hBF5OrgWl+OBwCBQVyBUfBwQorKZDZJlCR/Bt4G9oTZR2F/11
kSL9RKc3TqDK1Q1qm1ee3oPCGoJ0eca84Kv8nFxHvr4hDa4VpTYjSv5pQbSNpevfjJLZz0rynk8u
/naymmEJK67WHm3c91jKUKaCQkpUFov7S7tGi5964hG7TIG18/ssuMpayoWKeRz0TjPr2TndBxfm
vzEltEeWwh6Ij5Mme2QuxAO5HMCx94A019MHWGaBfohA/22paDywmWjdpldJCyPC72SxNcXPuHlW
OqMquM9YDjnFzPOFI6ENiOtCdcpbSYPM4cfxDz0mi2ay4DUuAoHe/xzeNpGH8jt1gkOS5XezJCNC
sTz4CZ03/CemiY1BCcPh0RNp6TQKY16o51/N0tgiJgoqDcXCunTpqqmHLkJjMrw/qy7c6rh4EJf/
qPXiOxe8AYpb1SPzBr4vL8cltpK5m/lYGLogRxJ+up+ESOKhXCsiiMA8HPmPrSfnqfSR0uoR5inz
R1I/JQNEfgf2/XeHpax5qzExbsayyzY20MfirbqP4TiYvsDNxhrMQqcA/JjTB0ALyC6SVIHASbsC
4HqmV8pvaQ862vVUQv7lC1mMo3CjzgESMwQLroVqg0ryNg6ZtFJ234UEQnWqLC5D8Y3uVlRtLLQm
1tGa+Fj13Ry7A/R2bvg9CU+3ffTHb1W/0iTdslhYyapT1eOMq+ZPCvDda/pTQUnfThiHfILd2Ueh
nxGn/CrLWeT3B+nUY24kAQwXHSWIrX5h0JS4wJlZ2tvmXRGcG3Gxd4JlCquCkl/L83a6k5KsRHvG
tNWxb+C5Uh70HPjaKByuVJLFEDe0rTF2eZYvqLr4iTXB9n59Go9wYZK1GFyHK+X/b2TII8o0VrXh
PAiSicrDaFaVE5EPXSJftMvQxvHdncWew/fRoPYMcftqgU+RgEDjt52oGNyA6hjzOhyAGF1u7UAr
BpjNUY7t4JCxUPODTLIqMdyzuS8AmruMN7QujjeMQ3EC1pjzmgUbUKpX5eMqkOh6LtvO/Pn7ficM
NPt6yBF6OM0k1+RfPahgkn22YSVatY5D5rau0yNDMVMHU47BVR0MM/k7Vta7ETLj1AuvV8OBmEtx
OQTjpatNJDgH0/TGktkwWjR2nNqNmCsPKA2Q+7GCxyXlF4MiAnAvfng5RDWmbU2eRmg+RdSO9cEF
D6pY5orYrhvh/XrZWsNgIk84IGYnI0YbMwxglT9gdZ9dO8L3+oNSGQa9/ejPx7DVV6LkLfKGJUZS
T5uurbb0ESG/DcR3vN3D6UQdEu7yCv4VaDfAYZbRbjbxCl+P+Dgv9syQycx9ftRI6OZxhmxCRzY5
PtM6GecKDJONtpzYW091Bf8ccWRp1DPbeYAke0liLxJbS0Od2CUt3qb3aEuvL9ZMkfo8Xdh5jh2/
g8sHf8cJzj5tBxU4iw0VkAeIm/d2c6Mj4MGUvzc58uO18uQM8KO50v3SUBMhd2l6hNK5dI5d9fq7
p4c2y/hI2z6V+1L4/svW1rRyHDp8tWUVIYSoReTSObfqS5X6+Er9IG0HYuj5MwWELpMX0HLFlach
EN2HVVI/7ST7yNFfd6UHg7r7KpYy2ruCuCelJu/VeW2hu3C7s+t3AO2rcyYOb22ijrGG/0GpiTvh
wU8t6yaMbhwL82OxWQ3IF2j0PNrbajgfaAL0LYNCXQJ6UBN3IEgRYf7RIJmmq+j+yvCKfUYLal2W
txMC+XfcA5hM0IVk97HuUdtYczXwA4FK2juKUKCKy7GC4InqXSmAuPHEbmpYtAC7YPuecRbtX6/t
//N8THzp37x6HrCDctqxJ14TDfwBuy0kV8i6bzGE0gF9E+AmQXR3rtHdPGcgaL9HoeQtcruZ42MU
sMYQDrHDbt8/TqOA8cprilWvGIAdiGtQBFaIQRJMKl1vEihRXHY7LaHKQ6b/3ieVZ6j/2rL5sBUM
oK4VPkR+qYOMUuMOx7PQJ0/PQ5A/Ecu971WF0QRKU5OMJA8toby0hFvMppXfnWdcayQd8oSzHzeY
iLXfPvm8A4uyEeaHMupDgZL1OyxmYyB72lmAfx5+RmmlNUj03pICA39W6m749qeBsNYWpP1NaqjS
GauqbDe9PdvRM19UnqxTZNPTn2Sq4WmgTlBxdVtu4qzrXBWLcWOvo+Xs2wB2UFiLrvq32HOagtjE
oM7wfRb0q1j9nTkkElA6u3D9zWxpdmqTraylbwYO531Wht1EOFeJDaERzGEHBqgsOFptD0qV6OpV
qbUvbggjoOLGKx/i80vd9bCYZQfW61Pxsxu+2c3ClOwzAq455xtoUpu/yVGudbOvwSHI+DTzj5IO
FxaUBX1fKyWnlBjpTh2Plln1hhnzELKdzhE0RMSFP/rnSdO/1Rgk1R0XDyR0qpfy3KqvdEnJkt0B
M2bnhMnFb1DM1sYQIPxBWQbydROnAVnA3cB5JjRPMZLw1TxQjaapg7U5q7rShad4F/irTmNFe4zA
FgY6qaNlSA4FkmUzD2TqG9cmHX0px3j04c9cNk82yovSvLZkkznF/Frzj+J3T6jO2rBqONFfpXje
IEAM1jTOO+mYq8KMwVzxGszX98VNqqnfzSNXXSNuoS4KpbMcC52Ky2FrTPtwYb+AKeRV1MqsLleC
p4YIrG7eMXuohiqOs+EYnDv0rsZ+WvbFbedNvCP0KQTR51LFHg+TsT5JRGKODqvh5BxLRLZZC6HK
OEB1JOtJaT3PhAWbrCKRwynodsivubNY2V71PnkR2GJlyDfM6y3NG6iBD1lTmmnqqfXu2pfxQE2O
X8EoaRxiwzg0Kpc0PA2ycXYan96Muq4pA2EjqKJqNzBfzVKtkkkrBbyZ13EUt5cSEBsrJ5Qz5O5o
WhaYl2eqAkD/Ped6dbkEEh5Zi199ew7+w6njsiSHu5r19W7xLyKJyBtTetxwvzepnPe4YQ7OR89L
wplUTtxfFbccvu2VfTqCiIfxrR9YmG0QfvJ9/sbO1JXqWWeJTSqjaW2WAnApHAhDK6wxthONHTw/
DPCV8PzauxnZFu4ciSgQbxt0+QazuBnZ8Bv/p0HiVLdRvBiVE0dgyu8jIEQucI5BiDjwDbUZrcAO
eivHLYq2ufA7JThV+IKNJ3E1GuN6P82I73keu0zEN6EXjud14OJIJTJGR2OX8tSeBixaWxuA2jpB
PciBzzhvh62uo4t+W8DJNbtlO2omEvVlOzpMpY4ZYJH05oXD2i2LWKvkFZZ++77DFp3g08IFnXtn
8Ir4H3Kt0pBWhDItfNFywhs7sqkOcOvmeBEN6hUoFqi0Vm6e3sFkXzQt3/Bu1FKL5Yec+PB6zx0E
DYx/s1vlMHD9KQgNcgf0L2kutuklveYVUWC7JkGSTb6UwBljI1Ax3FwyU8CZx63dS2DToicdF2eK
L3Dkrk418+U39kh3aU0rA+3ECaMkhmm2FETTpuh/Gl+OthCUGWEfg7KIoB0GqXKWZtVJFFgb1mne
RA+MHNoIcPAQlXg2GpvTzzfdtVs9TUYveBXUEdvg3Tumy+ZQ0uyoCJOPfLOfRT/7oWXrDt/3Rem6
n7AnS4TFK2b5BQzTMcSSqF4rJvciuaWV5tvZ7iASEd9I1Kz2db1KgGYRFPSSMOuUZTVrlcMRLpIP
RN6EpjbVi1O+P+5eJ7wmNy5nCtdYfSkTHpcyjjFquPY7m6WjpOFF/d3Etp3q4HrsBn8Viz8JzVHp
P8GaRa+z5Zd4aDUUyfiWelwkvOsx5vS1TKjDs0yHr6rSROVwgLKzqD8QG9kjhucQ1Tbv+Lcj5gCJ
DGwSmKvKDU/Vw58OD6Bh32oBkjJWORFXvVgp1q+cx4sxFJWuJ0YZX/WWPdraXNm30zcACO9sj5GV
4nSsKIdgv0PRWMtKdkaR/2z2vVe/AnfLBDErk99ThO1VRPikoAhxLpdvaygygRLSmqXEVmJXsGav
dtqltmqCOXFklraQXNYVLUGM48ZISazOYLRndx43/e/NQuDHeI1xoEBbPTcKeBgz2u4UlR6TwD1Q
1wAK0/LHurQatVriyNQ5OTpglXPACfVKj6B0w7Wf0x4qt8g7p0OOUZUOJlfK4ieZ/QZ0CPtW4hVv
vpHeQSKaddNQWI8D/sOhTAqEMpkvtR8YX4QVaZIBHe1GIawGzo+ERCsUARS5Wev9YaAK7vuBKDc/
XW/7txheqoj3bSoM5bHQrOsBMi2e4Yc/LCOU40BV0/0alOkBog8kdNinIx9S1Ga2xFuSXdYSC8kD
OSFwVmbG4hKU5jBE1fqjHW4MgB0wwiu4eTwNhtVpfP77tPThEf8SW4+vWYeSNFFWmzgfTS1JFOaq
Hnz1y2uTyz3uVrpuuoOt1e1dMQotds82v/2H1BxyoRx42InSsrS7P8KzR6V6d5eOUhue8ttIFgcm
/CBrjMLhqCUgXB2uuVdEX8HbA0HVIO3qWd95IchILXafJdN+NCgQQlPEbMclKbKwf/TQCL3TRJ3m
810XFwSwsxN4CR/6g9GPKn7nAADSLSAqrhIQNO8X8kAgWtJRWwHSO/H+4EIc7IS/nJD2Pxcl4kMp
Wj6EyPA8YtgQ8FYnPbW+AT5e3FPAuzm3qWV58ajw8r6weigRE+FWzHNuBE9oPX9a4P1wBTwRephE
4cHhPvXSTzfroonqhBj5N+zHwT6QFzw0cXOn6czJw8/w3JnSiueL9d9GFEKc2rksNrv1SXltQY7a
2rCiJX0lVzEpS5p649SPEL4uWMr0d0pYc8HhucpPHf/MHiq8QFrXULRPmyQQXAGghWm4HkR2Cxay
3weYdI0LaNUqhcJCSch/AqQ5hG6oc/8QWjb2xzOxPakAWpMYWvO9rh5OgIAtIPmoZM4dbaUfiH8u
UNMAg1LPal2K3JcVbkjoz/cVsalnilgz0cODuOL2PgCTvhN78P9GntRUQbAHeS4rh9TopmtoHpX7
S1CnHKOWo9vxJjYX+QNpRSSqnsP9irW++6+pyIo2Xh5cwFhkciBKXGWkoViNJyMmzI/lYkdTIARO
DDAM2OD/zRGGsYemHiL9U9kF6Ez1rqQmA0i1Ir9YkXQyI2n0IBWwMp0stH7gbqZjfV9tElUYhITP
BAuf2t1DDI7dR1sB3E2r2wMuI9rAxbTU1ua1JhbILRQrb1QFn6IZUSwqFdBaLYSgFhONpT0Xi7F+
uXW4KT9AqcsZ+qGm/ClDqGoOujZ3kjs6g02v0TyP/kHLzuY9B4fnSobWSioHqI1HcqxBLoI1ZiTY
AkzYVQM81N5TCp2ekNLlxbeHOOMrN8uweFQzpnmFQrxYhEwa3RELA+6hpUQoHRZDGaSA1ZX0SdDt
jzo3L9YQ3rHKyun3w/PN2zP8LDfY/4RpX5irlaFuXCgiLoP25WlXFGnxWX0bVxMxPqfLgLzlb9dz
wlsdNfO6O5F3a5kQD+pttbwVqLML0PDRBlIpyJVXVaUY9RJ87b8uMnS3CDk65q+EIbXpIICZBQxH
IQu86sg2gr01IudsavTN03GHsXRfd4HTb+WybFMydBolCEZ5SO5bocDI7pFAFSTp7QehRrOk1ABx
+Vh0YNaMbsuy6ptFJtLtYi4yh80cZvVXmy0mMwDhH2f+0aBx8wyOsDBgbLaPWKWq/1h6OTIgObUQ
sKqdm6zQDfJWn3iGfnsSr7RiivDRRQgHoIfghWkjYZikCsZ0BoCmcvRLDVEilQvhj2hTSY1wob3f
pJ4KUgRaFpDaDa9uT+TB5ztmRqXUy0tVhzRSEdZtJzJ0vDMGF4tWkt1aLxEjmaQ2zXvnRB0olNeA
xx1IVVrhJH07Pj6m1KV6fzJeBG/xrQrEzFMN1djz4dwsdKICPyPbwg8MwREjZtfHwVYu0o7CSlJt
oaj1HaPLIKZBNBpV0dyRfyneMQousnyAbuZhESBVGN/T1M6t/uQ0cHR/aQUizzUqx5Rd9H5w1dOS
ZB3wjAL7vExMjoXTHAiKmC52Oeb/XVznVT+c4RQARcwUm/U6n0L5kPUFR1uHT4/TDmuAeMC7aX9z
oks0Z1F8VEeVjOooGUCjPZDSricTtbNMVx6r8bzfOK55qbWC2SX4ilD+ullgT/hBAoKXp1n4g9N9
KFZJt/bNp65mAVV3LzaL7M2I0Mn5phA+mWz6NEwBjBprH+VzQX+6YDdMyibqBC8fH91gGOP6rSIK
6Kh7rERalcL4jK0jKzK5+qTu8xzerDGpucXH2S1mbccYK7HIby7HnYbybe3w6EGwHWlUjzvb4pE3
mxYo2HkAEZz1LNitH9J5arwoe5DgvyKmfuVQTZccUbaVk7MD/Z6NpDTx75sFHkNd1UIs1/W0Yh2n
uEOo0cSpdBd/o85G4V7ybQarzc40DK8zGJ3KOmo/E2/066GNFCnEds/lOsN07TsdGLC3Mndi/jyz
ug9g7qQQQQ4tOhVQgTX3DzsjjAzWPmmMsAeC+KTrbHDVnxyqOUMfMqEkneS0zVoTab4o2yBtUMg7
TcgHXFw3Tul0KlTAk+p4R39QtSAOz6P1xA1zizvDFyLz1NmMAXrRpObZA8yh8yAJOrN73JRBBk24
qCULku0oMeSgHlFhWrZmlBn3WkbUkZWGCTmnMAdI8cyaXKHzFFt7F5e0yQf5iKlHnq6AfnGL2nNe
NIKDs8fBkDLoLoOnbz5CrKhZsiVRvrvowhJwOw4kHF8O0fOu6dcYS9e/bJV3xLCENUImllGMeM7c
0tZIUqWdx83Koz/waOhQNZ5qObQJ1hc9u6REfYBfl14TNrk4nMekCLpt8wDfaBIJ3FACUNUPpDEj
zNl92eAYJXTnsKuwR3p0x+zzUp64B02MnuFlsjQdkaTLKTZhj0ZT2e7AYYtypY0ECsfRCEA163oE
P/FdvMHzsp5D3V+5ZbwAeY7dxzp1Q3iXzEdL/Jm6W+ZKkYlH1r/5VVKSs+rvAcsjz/hF7oNDsRgp
cVx3JJfEJ5rdBpJ2UTIz8HfNi98vxfZVdV83RqwkxXjtcIg/YL2O/APK9dbffs7UMnFSIyv+aW+O
bNlaje0g/1+pp/HotQdozeC0e2drRSJCdj5i4b3J8ESONBvVeXs/9NjVLRgPm9/6xs8xG8TZJQR4
opSZUW1JcwQpTtAuHT6yvGHpgibWH91aGfEW028kR9ad97honvdaFZKEfRSajP5F9c9ETW/e5Tch
lJLs61Qcp3hqIW2frNXosgqMRNxlUJJHnS95P5QcNKWjqEqv6dICJ0PLXTjKRjuk8G7SbtByy1tJ
lm3A4ftvxGZ9eu8Nvmb9Dmi+pWocGuE4moUolpx+6KawPM92SJuW+RSQoMGCpFTp3pfY7qAAs3nE
x3MJbQ9dOwlc3qv96RXEcD+QEamJE8OVKkMdMAihvDhtpnaqem2vAaBFfxBQisTyvDDHfKWz6lww
CHUUgsl8JkBx+JIM32luF8QJlJ3KgSck39Jew9f/+LBgOYAjZrq8WllC+SSL/nCAL8TuV3Pt2uaf
Un5FzXSXb8h4jgfe9gDImE7KbGPDkRCUBHJFwdlBxYAYJG54mjxbsHLISEfkgD4pcpy67MclylgG
JUBVXnb8+nk2yHXr/A93QrOUHnS2A0jMgVVsweEQ0Gm/swiRCj2qMAz46Af8iLeZCH3P5C62oVhu
0FaQ8jH0ZQgpBXLHvvFDOWs9jbRtl+9bxoSFBadEf6sN/wKy8d0MUCzcb/gDyYyFaeB6qknFQXPo
1EDRnDkPHdKqAEVdu11A9lIvK5Qroo1xrq2z2tFdKVp8fbRVRkeUvufDP+aw2WqPFpE691iLy30B
44Dp9ahJw2waGPkANCV9ad05o6z22eschIf5TYspaGPmJBkwuy0f9Ls9Ad5JWRZ4qkAPMV6lE2Dx
KEU00zG9fXSyM0XBjTMRTduurcDwyRPZP8mxSVkxaHLOlLzRrI9yuQygltsfHWnWvjOv1ZN2xdax
+rp507dUOf9jehxrMAdUoz6mU3sJokKZnzcn5bOhdJxWs765mbaFfvbFuiUIto02bXAMtuUdzq5c
5Y0dmqZ9s6tQwqxy9nb8MO0uThkXOC4YjxcAZpwHB6tJvMPEvnyt0mZOW4U8ikOOx0niD6HyPkaq
80eTdYwNoCuvzmwWG064Dp4A5ALK/sUZUOQesH5nYPkDNfTkWZ4QMNlAtqbCjYxtyt9hD6K7WJLC
TAU4st/+ZhDwIP9qELNLW0WxPcZHOdR5kByx4k32r0QL2cy6iX5Mwvm0LcNCheRXahW7nw+Krp9C
dVXUmyW1m/UybFmLEApFUnHGNVJApdPhbbImj/eDLf5PtkIrQ7T1JExbARQizPfntAEdHx7Zrbs3
Hfk5xnYNUi+2cE4hByLZfBlVWWB5WJqx+2xGHCXgmCWCk5biUNgZ2nOyVQEMMeiyZfVJf5lmewEN
eazIHaee2izciLrjL3U7RpGzu9QpS1o8OD5L0EUR7AJUA9CO4JYSxIaaRE1SoQCzn7buR9Pqoccf
yqpkfZg52bdO4KUDW3bPBBAKBRJ+GfUl2FujZWWNegeLEL/ClwEoYBiTLfH9U5hpurTNHnQpqTG+
xPlQ+xpgU3Nl0UE6JkJCLA55keAIeeQxpQ8uyoBzf1eCHZX/SFv9f5dIdY87M1xazIkneCfZWhkC
UIhEdMBWndGHvFWB85jG7dh3sZGd89HdqiSk68uHE0PONPhMqmFqQGVj1SGgWIjgUpnppkj6zqrv
DR0A2qA6xKYtEaoTyLBFRq8duYd1qdWMuNI2I87tULW+/0ztmJMGjS3wF5QLq0/pZPdW6mx9NxnP
kkBTU2a9L0LKMXN05NQcyYK46S6kJBBQuuwDWEP63FMakFm7XS9aGM809oco4dlconWeWB+oiAiq
APMVUp5dBv3sWpC/DRVPhjz5udaMhHEGk8YjkcgK7MemhkDKcIAqLJeqPDxyQ4JMSQbIyrPaLwbQ
CH/9vdEblApBbQ4d/sIZ9cdMKEb33Zd2FSbAlv2UiXluLLEq5jRtZeBNlDHwfEbM28gkNPQYxcaY
VUHBaPjBdEUKT46qd72KM/0ES+ATxTnNZwEOTge5dZOfvne0zFjml45rLE07gXep2dbMSXxjsI2o
UCI8PYtGKlOmnDGs2eCYcgoWD8X8JyGjVhkXl0tf9V008uLdBJpcUU1hUCVcBWjNk8+359otmUyM
kkX35u2J49iIHTneZWuC7+gNAx23nS/9qT30BjGSkodj4ENxT5plB4lMwBpySb4m/B3Dm5TUDoLy
gISF10KtUxqkYFykcQtUoY7OnpOdGBw+bQ1euODFGkzX50doCtYPBPk2rr8cAZJfHzNqXTUQoRaQ
N3W+BWMZbzuPvDIjoRaiN/H563iussu4/lASsRM9UwQgfTXFdQ24z91WpBjVSTkFFPkEi4cbd/F8
xKnrdMT9WVM5ol+ISUqy3NJ/j8dlfvU+WKOgdQJAcRFuRQ8JK0MCrw3CywrlT1QHwRxGStr78sIK
9gQaKxKkBPaZwpdFFeif/ZEwBONnjeY3tJJdQxg5gbjaLRGkBANrHAVgXGIX+68v2AQWJrlk4YMU
3IZGt4aanR0sRufQ4Ogft6cMDy2xNz/zN3tDVFCCS/MKEorl7jNv6Ax/KBZjoNAJmtQrBW2sOHgK
p6JQuK1auQdiLFKOiNhq3DTL3+JjOa9fBFsT1xPBFI4oWrkN4U7sS1VIjbkfn5yTaq1GEW0WEOju
kzlrOX5VyrRzZYVtP4M6ASZ2dYvdeTQehOfeuRbiITkI/jTMbsVeyOQcV5SqOBkbTRGrlXzGTSWT
PmQS6vPNfRKPck1FVwSTz1kpsmpwbeoPJXRX1/6D9t5UgmZCMr6iq05s1R04Bf9V5rmNyPLkPec7
dBri/a92seCarspi0EcqbyH8k8OG81Z5wgelQIxLSbXR8zS7PWkil0OZyLmMXowq3BTE3aswoVPD
sf5Jb5p10K0zfeAQ4gzSJqrIcyzu5uP0ItZzroJ2M9hR+wad+tFTm7HPpc87IlyoC7X4NI60BEUk
RXgDIX6IB0BrW2MMG9rG1yd2jL5Ay8FD+qvx94REiY5ZKc6cCMjNLwy28QRTF173kEQea2S7KgA8
ZxiIA86Yjg7+VSPntgD6MaVivf4x3e+MdfEhz23M0kiYFEsBeokEoQU12xeZyNPJQ/4c68aazVoP
HOXzgvYBCrgB0JRmih1UZDiIM2BKJE9Y610UUrFKQupayvCbp4GMX9Nnmx31FjhE+jdgv2q22+33
eUy7dM5us0YzTho7Ykvl7OC/qKhofBjuH/BR0Vvclj7B1ku4z8enn6EJ3X7u99l3FaD6ESJUSey7
McrC1nvQ8ehdlDAugGC0TrULCUf9GkGWEZ6nV7v/yDtie74jx5Wb3KgeSwlLOWtivLVd/z6bdNAw
ZI63/Ij+a8biNHFSyJN1uLB8T/jALWZKmn/QeACbVFkCkH3KA52IXYODgxEebzZG6iJTqF+j+AL9
D0F7qlobGywiUJdh3opqg5Q8wja0wU4soHrRK8ZsPeTwdFxa+g+ALi3+zT1A7LZ6gPJP8oKIscP3
BA4wZqgE3NpKPO/IgW1h2PCPFlPr3J0ecJE0CJw123lhd/vpVdXDQoCLbazYpyzTuSXy5yLXVgi3
dkSBRXe4L2Eg2s/rzirCFFn1hKqZNBsprib2/YaMBvWi29swH8QN9QXg1oUB7tXW51aXFjyXENsT
I2PgWLost3T1k0FqMohQ/qyO+1EXRtKfpDYQ0v+FJb1OBjtVA2yqPViCuk8sfivC61EpC6eXNJ4L
ahWh3cGyerY/OVfZKFpwxEclYusBmw12YQvlj/YBJ/rCXqpcnGMtjdOyKCVb12CeZS6D8mPeqnbC
so6hyYeNexUleCZJCMs4c4sI/Q/Bi48akH01eGDXzIydGhXjT+vXTGG2w7f+MON0OCPjH11fCXt9
m1CCye0GE656qXkItkYGR8RnvOjY0/n1kBLudetR0RLKN7vw87dvKfoj7oKdsoxdAq5kGqzRh3rH
jRFjMgbzrFOxVSPd/WaBYQA/CgZ8IxbFH4DwS5J8W1esmr6JvuOcUv1PfMBopshbPBF84Bk+hLch
dranXFo5QcXvCeS43ZpEIIH4bsy3JVBBLvNDtjPZMo+vpx5nB653ufAq14VpOmB7HmruAVUObdwB
LUTyL9kXOOBUU2eKoZh4ATeNvedFCFY1uPrCjp2HNdK4wWbiGyQktzzo+RJPIzz5H43e9g/uXhe0
r+p0K0+nt2DGfxk/SIrt55F+FFszrWEkSgpBVsG3cjjqNd0MRFGI4HDosJ7xjLzLVJHAVrcRbQ7M
xR5TNd9WCJK3dm+bKobu8gEgkicF72fPwFJUhuBlj8MqCBdxXbYh9yCXnVY2bRCQ8sb/PCDohs0J
DsjMfn0RE31ci3iJ5hmMYymOPgy3FUsq9QIxSeeNu8U6V9kbnh0GFjZdYySZIAyan9tCS0Gpl1Kn
+jzNG8zPnQmvcp8oA8ZK/KavnyiQMai5BV1RFt/0v7Wrwnb9M3fLXRdG5Gj4V3nrosBpNdmPDpXP
bpoB34HpKRRy/XuwJdx7Xc5jmkrC4PAx5tpHuvMW7tOdFYsCX33WrOKCqZjUUS4MQGja53ss52wH
HhvcOIcM1UDY9wRlctO2yebQyAIy2dWO8LqPbVFhG9UwI8+jXAYB6ovZ//XI/RQ0tEugAQGHQSF/
ucCg7tGcdWd35T+uIOy/ytStagEjbTX8Otl6OyJOjYvRAPuUjz72TJA4yp78TwkVyIxfdUY+nDaM
/438DHGGSAGNcLOe1jj38YmKqRLSO12aUA7+NK2/J8l41C/Bk02GaeC5lk3Z0kX9sVUnN1wpY2Fw
zIxpFVUIbobzSRW1lQuTH2SPk4IsDnw5vbs/ho6NC1DgRhmzb/dLe4m0AZ1+JAAr007FS4Jzk9NN
UjaPyTpkWkNOPRwRMcWCjgTs0MDFYHF3p2+mej8lZr+PZC9bXeWwQf6tMulfn43HgRZMM8HkBbpL
2Iq2pLze1p41ispnwfCT4/tAsC/and8K4nspEv+IZmUvPn+zAtLN5VMNJKBEea64ezowC81IGvBN
ehYjYdEE70K+xGG9pREO8hlwxFCjn8y6ntcVYSKFDKrrWJOiD8MRr0eLNxYsYhQlMAFmnxJjWd4h
PZmXrw5IUz1BsaK1wkMHly/DIFJJi0Xb85unOGP9y9za/p2F4zNMJdE0Fncn/KHJXrrq0qLZlZrS
prag8yt8iZIZQCUBMz6Cu/O/32sZsAvg4gqbDRNRhXCjhrwkUSvq9isS0ipOk8cnWYC7vYjHuzwJ
qDJEo0jkN+PIegbgh/BkiwnNVPHRJF2HuKsxnWcxTWcyvb0C/vxso4IefrC2J7RyxLX1YTwfqcY8
x0EEkzRDtGSS459dE/5/pCY5s/MRbIb3Uwv+a3fTLkZbqPQe0vZfGmgQSc0gkZevgFUrgMyZQx+G
u2bAfg8Q0vj4k/tiBpnsufsK9gZs5aaZ2M2nk/+xGgo2YR1hkGs71Uz0qG7+B6lTb87MaM7uNioh
0BMpDI6npnXR0cKwSmOibo5uR3mdD5jKnWN27XhNr40nlEUJrnbWDdaGGVJ8Zv80lCKu8cO71acQ
p4blo7JrkRstOUiIpg1ptXea6JlYIbOoZYW1W3XaSN9v//mptu1+eSbdyNd8gv3zILiNr8VtvqK6
aWazN3XA9iAdrOdtOURyVL/f3JndGiHBaJY7/+ZZQ3OAMWTzDTLtYJ15ibYx2IH26x4J89VOlLTs
kO/8vGvTNKhpGXk1pHRItodOnU/YdHcEHmNJsd7zCA5xIPeaL/ektUE6NnfC1pngsTDzm8Iov84s
kNFfK7w2fSZrF0yy8AtHqr7DgSloxQvzKm4o7VJJpo2nkm6HMz7tm6PGkgTWG3C611YqTyLXGnKf
Mc0dS1vx8gc9lKVtu0ma0io12IRPErFaa3lxeHlWUt4R8HAb1zsZ8SnMV/hfYMho6YlciuyKM0+g
F0kJSKxHmGWD2xB7NQXFL2C5SqQPWY+Zv+ltBa5wM6RFRPha6DIJoq302Gb2q/s+NtsAZA9W84ZJ
32FvXv3qko2jiL6AERbGx9AkAzpIzhRR3N/OUtHxzwNpBiK2JST7PqGUNNjtfypJIJd8sVD3191T
TuQN6tRHnLbu+n3ceUeNX/EPUnACJnguxvIxfp8rUUtSPSFR8mHMpUcI95Nf0RCPLU4c2FThRd1Q
fBxrdr1Dw8fAAdFC42fLYr3IqWzmnP4D9nvVFzKnuJwwyyq58qzkH3G99C007QgDJSl7cLWamAK7
iPcMRLErTGFoBsJWNr0DzBX7fPQds07rj6XsO1vBG5aQ59MhVfLJVVy2vVUVltR0QtWmUxts54ES
f9LQ37rinX+Nkm+G5KDRwTS6k90qsUSwZi3w0dHSUnV/ekBh0wNuznQZaTQfpSr/AdZJS9TH9Mlp
3ch6TAITPmH5f0iR1+uAv3iPA9fE107ihlRE7yUfFaNTExna1jftA7pHhmTioXSyE7cxlhxdzGOC
fMU0kuR+vy3L6DwUAF1GZ9AdfR8H7Kwcn9Vq4/ODgoNioeUat6p26hKpQQYxgFNM+AlLVeV/vkqq
+xIyy6Xm4SCfi/b6DJjNzxWhWmq7uvK1i9H9kHHTVpEJxChFDgcUDcPARWjChf6u49egxhs8jaw1
qx0J+34v8Kn2WEouGA63ez7GxEh+1IqBTWK7ZFOB0/Cy0uDCDAeX3VlPG1E03/g7nvNegyP9Pwnp
yx3MgIYrz14gByLB4oG1SY/HVNgTsBWp8Kgfd7+f0CIXGDV2Thcm6075jCBjWvHC8CiCmrLZzgiO
kZ09PRzmlwWd60rG3tiTJa+9pJMqtqLgKNioAXNRuT01LiP3g7i64+WW72lMpT3vsVVJsqLU9Bva
AB4HrhtJrPTfPMOr468SlW795LzdpU06+AnoTrcNPM128mB5C91hDYFIyx+fXup6wpKjGAXhNIKw
QbxTEKPJuvIqG8j6pFSzYKFS3sg9HTsU0mUhlIlgKXbTqoXehgv2L1BRs4vH78CYHD7Re/++6uEK
+eUwa+4HAEnqznDsOHFU5rZ/9naiYzVFpwa5V4xHPcrb69AVLttk8QJPRCvPB8YLAobrgfuNwzbW
S1CXQLW7sWJeR1APz9fr+Tv0s3XeKAp0RHp6s0XV8PaRiz1wrEr+Aa344zFpdrx1qhaufyrMQfbp
tF9gBPJoP5PD2UAInNXRYw53bOZTMkRuenia23BvuvOLQuPMczzVT2MP7XKMvbJBBhK+6RfQ/Jon
FknS1Vq+uOcHZ14s6La6jJrcnb/Wx9qTqRit0Ar363wIeeKgsdMLHQfV3oxedqXzjcvyy60MQUMD
/xt3bEzo6npYh2x8r8SBR8Gw1DGaBOrfQMGN7noWmtES4Rt7+LDKxBo40ZfD/GNZVTlUsOnYA97H
vKMO/lVAp8m5DSt77TL595vkJoiCJZLKIc4o4EDKH0O0wnzqs+JUWSF56jWprcq/lhP+pVgbQnLp
/dVYXpDc9Lh7CXnK31IW16xqJRfxyS01VDHS5KimNZGvZiFXDfZFCXKFzCTdzNLQu1S7d6KEp51p
Wh/WModveH24RXjBmT+z3xHfLy21REz83vM+z55EYomIrwZOG36VrVOdh2n12/mCR5xpyOhkNHIt
TIiHnXetScdJ7KzwzWbzZvTcUU4XJCpRXCq78YgZ6JkP8TvH/bM+LYO74FXb2Ps82kmREHVRuIjj
+jlXpiIQOQocz8CflkUZA/NXGEmogLTiga2oEXGYAQLCIgCnhPY8HNvPVwBqt8bK7EFRx1vuQ1M1
2ykvYvHI/KJCBiY8XI+vJOesRKUAlsDdFv1WJXDbGB4Fx6/mSpoov+KKLbLNpLJ8+bkhmTR0nI1B
il86IHRoLfvUbKH2+Pp+31jwv1kZlhsWgpjK3UkSZGuHO+dS26zwXomziofJybiB1R1ExTPh8+bF
kskNrXKogP2wRghp9jNH5M6WHoZ/6SubPCLwGMUb2tK+/99I3EodrhaK85xfTcJlhL9SHe9l53lp
/et2v52uKhba1aeW/zYZROy7TIHt9V3HM6+4k/fLyjvzEdvRcCQ6vlkIPdXrLKk2EEj5r3v1GUjh
vQyrS77K7swrUw+dn344W+qtBx7EFOcdx0oXuBJvRLCw7s1oMtq8zkAtbKgza/p21+M92TAEboMP
3Yqdn3ya2yl0GLGarNmiIL/H5heRI15OlifZv1CQZZlArxZDX+jUDwnjiAg2IxO4hO0dV4SIeEFf
wWnU0mQQ9LWYv3Rb5oZa/ngbu3ma/+x8HRm3k9X0GP+g+43XxF8odqQuGyVa7K9YB7sQyxlmv+nD
NIN9oTZVID8cjqhwy8c70n9TzmongsM0Er90pQY9mzPRQYJc2xDxM6QoP3++V3weRZXz2Oxn1urt
4Wz47Oj8eeTlPgwda/4D69GddC/GvuNUcw74FdqMPuctzRVSry2ufODdlP+VmRrSZGvk7KxS2jCQ
jInOPuEgA/hNCUU+1PtfDcBgMUgiIpi2tX+CxCbcgNK56wjbiqlS2k3x6VVvC9HdcDiVZgRS1rsB
6u0/AUj63CON8QIAtlpc1/gv27ZrtRzb0jt1KT7Mz/ZNH6URduL2AgIJQQNPTZQdKj+/mOPfKdUZ
UhupCic95Rw4uGT+DILy10Fn17kTnKSC3DSYwSoXMJ+hjYrYEVXqHB/DSvXlBJzfSAa5DalI4XjQ
0HsttosTTFRLo0tY/4rOh+R/CzeADcM8pzSRHPeRfPUlHGKB7FsTsUCr4yeMyiLXeKxmPJIPA3s9
BLn+qSE5ZTaYzdFJNjDPDSAO8WQSdpD9vpQBWKgDV5PDblOo2gL4AeMXpMfHtVXBW0YHdny8mO6Q
WP36136SUbnR0jEjKOqWnRSlEAgQBcOX8muDJTBndT4GcmgPHkMnI4PIKsaRaxPi4yLWjz3WsPQq
+DUQteDfuFDJKfaxK72KKqDR6IAKaBvXoCN+4gB7Nb1ezzyLDB+ZuJDdFrMGvTYxERND6GOOa8LQ
QQbF6z/FKPGyhkMDLaY3jgrdAZiDAIZv9BjH4pLs/Pslyoefp+DJM6LSG6To2USz/PwoeK1FOcCO
EwKfJmQZ3XhCiK2Y1GZnOYDG+aYWIJpU5D4PQsR/HfYh6vBdHalQTEin9tGV2Dz9JKQVyy8OSJaO
8u1NTeffxO1K0Gd+Wu+bZaX9+fQ6YnCt8fiJc+snpsKG48vPig743m1VnjWHQ1W6WnsyJ25gZPzl
SAIjsLdo22+4k5xi3O97rcHxlLIANsdzVL/ttgf8BwD5W6V8GuonAXKWqi0Cd1QCbfzVd4i8M5P0
TOJlMWa2grHfgjSG0Ukm3tHXgApW32FFUC+QGf1HsOB1jb2JeYw7/K6VCl0frpz7fQsp7CiQA2MT
IOgf/wc8eeGlo+AAsv9L1Ol9e0js9h7WVxvnDEOSRJw/WVlA2orw1h270q9/WYC92+IKNID/jfPo
vzo0cBngU+COvYnMpt6liZkX+Dz4x7anJEwkbMnAgof4iqgQjRy6Nf5IZnm+MNkzH6lD5KhuTuaJ
Wr1+a5dpgf+GKI6S0zLRFlYKnaTy3ZQwD9q25IFoK6Fcr0wAjA51HKma+2wqAuKNQwEV/6Bn6v1w
U/ceJ/lXEyWO1U8BGZ6ovEaE68GjvAsWqf2K8/xV2YyqcHG2ukK4iegb698p9Kn6qdbrmELLdBca
BzIA0oZJWAxkpn/MKnRoBQhQ8kJG24LEfJZSLSeQ5JnK935KT3+kUw0lcwlxTi8ywhQDj+UJ81o3
d1+wHZCNKdwfPipP8oH1jshHbJGwdESBUov+VvbNxLGGN0deGjRxIJWEbl8rknJoOJzrpefyAGbK
msw5DZKNaQFMuE8fnUC2paw1isTgnSxDQZDKyq6QdxZnaHdWDswL5tuHgvgUUbH16CdGWOuUqi1f
9gCHXV7FU3S9wWbTRvx9GwRfdHd4ISoBU6XHF3EofigypZM6Zlx/49kymn+SjGcqpUxN7ksksFzL
wikwMe4oIniXl6nAl6oRSYtI4eoXiR1yBYxTxIyute8o2k9jVFSqWR2wbcBmUWVwHpPp6Id58+Tx
aBcvB3wAEWQagYB/WxwbP54Js7QwBc43ks+MoG9OAE4whc5wEic75/FsAl9p15UInob/TGJKeHA9
dAUZung9Vpz9RXy/M+fTs8vsDOColynLVCTUhZNvWRHfEKwRqylSySLejy7rVrcdEaTSsPRkH2DI
brKT/QCiofwZtZCexfOo+PWPyzbvsJtV+4eC5zooJmrVLHe7OtG1MsrvdtsxolQvpYSVcElvIgsy
8+tiXn7J/nEX1oMaCz2drMzQar9u24GMQ0k9vCOjY7zTrvbO9vRlEWpVV6GvsKGMFBVWfRg3GNGU
gj399Jyhx3VrnWhWyB4o19GlsVjdU/QUF1+XoKmoXhGyKI4VfXh3NtjfYvZi81nnvQrc+PUDMZNb
/n2X2BPCXtJptsP8UIgciOGQxt9/21/WJ32Yyzbil20xMZ9H8BnJRTZVRGcyxO4go4CWipDMonRv
qUbM4lqJdgCrBKSU6tCcS4jtwb0M3vQt31S8kZx7//JuH4i8qzxjHbdSHKrkCh01Q3Z+k43dNppV
puGDSPAQLb9iQ5WIv17v2kTzCKJHjm0jaBtJGjHCPKRjkxZl20xCAm1qAOI4L/572ZQ0S7+rotcW
C+Wj1nykF1jHwFDCRE/nc6A3BgE0lC9liOouvarFLYZWUdCqjM9Xo4ybQt6kUJjXNf8fNsE3cK9F
F3YHnTq5xQjDUyhCDtr7YsTpXWeO1eGy0qjbNYEP03v0qFgExV+Zfi8UJSyzuV27ik4fWlKlUQFJ
ELVUWndhFA+HGv0wFbjRK90C8i8tkU2rcz5SZDHzZkSp/W5hJ0UaAiHurBQUbfYpyKO5KoEB/9oq
WRxs592qyhCrJTHCmhWJ9q83PBIuMOwmx9GzEvnpcC8E7eyDu/TMnkjskDE6f5p3yAOkrb+6apuu
xm4bpxAo1khpaTcQh5uXVpC4lI1KIuSJCS+hQX3AoDyRNciVg1kUQ50QMCnXRgP4C8X5kXaoNz6Z
b4iYKS8rmF++Hy07HG34YDV1fhAd58ndULACdgg4w0uWh23doKGN73Vi4Y+zKCjYvAvEMkBD3+O1
caHR9cKgfc11R9Fi2Wx/lYz9DhoVha/XCjolW32ruYXV4qWMCndvzvIl35Ze7Agmq+egJblItY55
n75a44eovt6U4buc3yygIrxb389Vwe8OyIUSdEwlG/qbmVcu6iFId7TN7kdDhUn4L8E5zLBN9nbn
XutzMvhoq0XqQ3Eqpx+P9o/RoUh+OE6+rI6i1XI6wvp1cb/VT1WBMDMrDiN/qmfK3V6gqgmg8cMD
xYm646xOEfdTnNg5hbx7g1XIVzjhoUO5vzCUQqf9TsG19ixJPHYb788RPpeArNUAmoT31t5/slIv
qlDNL8zNwmT+nNmw3zLSEeiVWriCoWtQuWNBIVHfeJQ9VGsCUjFyyg4lBWCh3Q4KaZRTQMvhPgbK
bb+fFacR66QHqiuT7feKIWS4W8Q/eeKA6G018CBBHS4AawWf/jzV8t7DUs7YXrfPI6xiLekppeo/
mWv8dyUyW2QaMivK3XQWiBc8pEqIukk2f5ObRNCrS5eYpoj3zPTRiPjjboX5ZgIGRagCU0nidsH+
yO4vzk+rfDf5NQU/rrgoZKteZMdpBV1lOWD3aSs94g2V9zbbyC1z2sbAVUVaWecZW3B/dDOortsx
gv57feeqXuOllTzXCEdNUooy6iOI49ZPjEIYiGvsLjoL+GlT5CSaOmInYLgHw5oaLK73kFPaLh+3
SG9XfoNroU1FXk/omc3L7s1FpdWWPzNH4Y+FIUbV+fbIxZz8Z/POUB2cWgABpCZu5DPJ8D91Oumb
r1BhHhYPUrtFIHoa0wWz+LVSxmP/t0xfRtyyB4gNw1mBHSz5BZc2FOLI6VOBIy8HTeTwJvfSgTK/
E30TI4Mq0Z5tEbw/6lH/yozU/v1fkhCoHHn/HCMW1skdACaQc1uO7xPGhwc3g4J4r1keX2HyrZtW
L7OGWKw9sc6JIS7a2H1iWr+8jA/9vKgeJQotBbMI3cT/CjRsK0nKxdNL8xYtQWRlnzvWCShkUq2G
8wnASdWgN6AtEQ7iTQuVqOoQFPiSC0AQ5WQxXzUpd4LD2tZN05yR0AmQ89sAkYucswLENOBR0WLY
6rXj2SW0cyCVFgDXfkccK2ekmdAW0GRNwjwbheHb/8q4xWCjdLya+ibXjQTjVzYe/lmG1Unc/8eD
JepNYlmq2rISbCy9488Vo6oj6YY8Sfu+wYLrMxhD+jGQgi1DYQReWjEUhG5xUz9JXUd2wIgn3y3x
iWiUaBxFLueb9nPlGHGMANThYf/EMuQItBZncUZQKOeJh8d3Xr/xEsFjoMItGVGfxfRGkYLmolWA
pCZYUtPnU2UCfGSiMPmrMWirPw+SE+Jt718Ums6Ikq913yFQm/61m6vu4P3jZ7ptTveVIGnOhsar
FxwAThQBnHmM2sJlMyoM4TX3XJU8BUTKo42V6/83BFh4KK3DQ0wTtE80FCaXzNmDEWaKsfAMYyD4
kLZ84HH+nyFTKXR++tDDSep66RTEPcCamJqTY8wyDM61WDNWrtXUQaM5n2ItwKapuMIhrkurYAqa
wLZzwLO8i2wtiwOdBtPgNvC0z2ZB/7KJCj3/KqBFVakOEFzg03my2JArLOGQfR2k+7EiqDwfBs8O
mMWR8oWWlwWQqCQ4Ti4ESXD2OEwKFV+wxqT48BsCmwHhWiLl9xyERYpIB4OexZlMyzS42GGc1Sde
yMtmATyhEOUaNeujP0OiNGHesVK1EcFiea2LNGpN24Aqxd1iIWGkG6w04uhLMqS5kS3FWPcEwIG0
RHTbm0Mkr6CWKOtqHqb/z5rapKYyYMbZdV9uMQY0/lrIm5QaTA5PYYogGCU9WN3Z0ZEcUU32XQzY
UU+yc7fqkHLvB++e/YWAD0Payf5cnhX50dRpPQwaZ5ckS1qRXIqPGtCKXtdzATymFMuow8v9eqgX
H0qmAGBoA+EKAn1YrTEl/iedM/DVAvCqULhT2TGlTmarToqBS9l1moF2+1w/73R1qlWzaVgBt5Nb
+xLGl3+77ZQsT3yVK9gFz7aPPmO2tZ/GJB7jVO4vc2V+Icx5Bfyu/esWa1mt8ehO9571tiqT90D5
GbFas/i3pmOrAdI27QL7ZiFze1xBhQlbWGgVn+C4M34ly9wzswjbrMQDZIKZmyBYJR8mNod7TfV5
3fXSSH69bkgymnF4IFRgP6IY3BAs7gPDl4MLMgICwUhXzHop5SDZT+Kso2gSX9P6v7DJX/zc2xYH
XHZYxEnXKV2cHgx4dD3uRjslFPVMXpw9mRTt4NN7awXuOCX+qv0mdw40zDQB9DYgr8Fs2GBrBH2A
55YzMXhSKlu3qWPnKmOdwiNbMKccph8dSJ9XXYZAWP3c/Tf6Mu7omjYX8MpTTzyGYZ0p6HBQSxyO
8lbVQSjEbmqFJDAC+J8HL7aKGH0UxyljgPORLBQAXnpMhV2h+ot+LSt/ErirI0yEBC8NOKNU3U8b
5Igs2oU4tM3uo0F0YBphkUjNsu82ot++JeFM51/Ux2tQRrwjgIOV+/oWYs5YCZd8TbiGpjKaciBu
1kXc/82vfsCegoQAXxl721upnHBnhgTfySTKXYRUS1xbQxRut4T1+6sDv8RXpMmaw8lkgvv64R4t
2NwpkcYleOba4GfDyQyWfA2TKpy1pT/JKH6L1xJ8zZgstQsbF4n+1gbpOznUSx6gv+gSQt+yAEC/
RxpG0vB4xXEenga6nnOceT9I6u0Hg++4mAynok8OwkUDvNy8B73gqUrA+QK12gVJ5zkqPwz7u+Bv
sE3xnIwUxddgImd2b5M+DcNLe4gNBhHG+SnFTYsZg7NT+1xUMtbmnNj5sZv4pUNCvgZnTUycyBJt
QkfDdVjzjCIem+csH/MK1UeMCSOK2E2Q4N3aojQuT16jztVOFaSmyK8djJx34SBVswQWha1Gur/r
zCx29Mek8Av2+X+WEG8afxg1dIJ4rYRRnNU+bdfsBDjgqBmUekqO2vsu9iZWWVROY4EeeJJrI+Kj
jDU8/ph7AP5S1oJfWxOUN5Geg7I1RKwZjLjU7TqGTd9gEeyhBZZUx0GQ4z0ZUW8JHKVgwzX3x+f3
4XLGOTV7JEA8qFxw1wcOSy16xqAzus3b/LzM5YrbDSxuGLdedCWZiazAz4wpho60EC4PEeL9pyGQ
yF9UwAeernHQBk8IH/XQqFyjEZ2w1DAp73FywvInvnyuIpLF3w6Z7ndz1vxGlzNRioSBk+ljv4Px
6xhMgtVtxZ5AgLzd3xCXr0K46EstJANoUH3Q6Zme9FMdoveNpAb2y/J5+rzSFFPBlMxRD5MZ3n67
Ik8LBmUBBTp4wW3moZCUbdHk0YABBP8zEbLg18EAGlyNmohGOxrCtsmyA/VduqeS2TBal2/mEd0V
VOuXmGa6q5qAbJPVw5Qp/P0fuBQXom7x4lkcA4/FoEs7KrnNtrFn2e1SxvVWBp51is9ppj9GabQb
RmK7Dq9Owc6YqbOfbH8384znDd5VHrdx3dS1lh1f87BfGg+wfpEunbv9f4DV9K2s6BjuCw23rXeW
QzQ+VAMh2h+movPswL0wujI9sIUKm3LOHKncTJEdQ5DO4vayEMkNNjpxtPjRLrSxDlgD9pjrE4Bg
3jMeUG60Jl/l0Bb3jChJY6cBu3Y43Ol2mD4QDrkdQyz/LHUrfGjPlL3QCwu5etfAZO/HmxAhKzgM
U1LYFok8LM0Gg7ygSeac58RccM1FZCTI31lvM7kr0gez8OsyfHl0nMTZ/tnlA2pGYiJMYdcOFkjA
VkwU7fBmEgW1Bk7iTvQPa65z0GSzxkt1PfikfP0OyyoMq6TmUql+bFkHVmysb/uCeEFuEqNi9UHQ
cYRAPSES1r0aRrB0xVl1P2UJsyl8KOU7fYUnKFLfhEtBt00d/T3hPNJHXN+K170zk54ZIpqwMx22
sEsOInz7w0ZCUzuvqPxmyr7pmwRwewKqC8ofyP+797Ybd6b9LAOptMci9Waa7+/QzzUm9ClABd8B
oGr3OXxy+0Nty4WG+Ms2/c5CoQ/MiMiLv57Zio7n7/OQHnvnrcYH/fPm5X1fJCR/Hdtk8mhDkNnq
2Xbh2aMHUvoItVJIIF7yo+Icq2iyNZC+7x9g/knrWIfaC9gixllisOq/vGJgpB3LpClI/gooMGJO
BSiHfUNRkBW9mtifAdehsnv5E+M7xos8IKwxgVOvjuAPRLLIFCAqPv5TdIlWunTZPykiaJ5NG9Ts
pn4/UTZd3Rlokc9OXHQhese82hQRqnM4yUutRGzQlfds41AQWeGXKWRY+B7M/dTAH+VCsf5FELlW
F7hvQ2BwromaFDMVMrsPLXGHKPg0iKhEFJ3v1E+xcEuzibAxjtwpDRdkqV5JMgoxlJ6ftdbmlS4R
aqUwLXg5NNY5L/IFcb/tKcmiD5FiUVsF3rc9Cx6sJJIzw7lCBYGEAMRdWlfNS27zf3LT7bvkIYrl
9EdWQ9ZHTs3N8VeetpHYgtSzlxjIo9lyIRzjB9w/EzmQXeHqU+dDX3aIAIwC+VeNXQZwAxtMI+1i
wZRHFWKLm+BVHJyuBsgaXLAmgJRS2tVs17YeCePcoJs96i+uun3PPevYRN10F+O/R+TkT0atJah5
XARt0/udMnTqVEhmrBSe5Npl+vr0KAta526fbQxqYsntLm5PUK1EbdOzUOGyyRDqkW+Zl1qE/sxz
mtZ1p6LcXeQB4YpdM846nHU9T3Dum9pBXcANIMzgt31kMbbmF8CCz3MwoF//sD4Jjxs0c4GTZJKV
m9gYGKlIj02apHhsHtakJwHVAF/vLOLJLdA1Yi63qCYZfPysA7M47P2NR3qUkQ7d3qTYv28PQ/Xf
LgiTFwOXK6p/ANIfbDZDLd6LjyIgOJj88ZV60B+1LVZmA5zR6Ay1T87BIDUrgnC4e2R6ykpQlnRi
1TCID5nIbSVzYoAGiWmYLv0u+JqvUcVp8SFH+s/6oJheCzzydw633ke5Rg9eYVwS5AbH6WQEmxok
/2RORbzlk8mQuOWJdiWb8jjqfP+E/5wDS4oO6drrPWSr6y4nQEyQo8hhEOyCevHXVpi5qjtk18gb
WHV0j3Wdb4I0Oo8w+rqlV0FXNHfyZOXTCOOUqq7uyIwgelOcJYeSR5sQgi3GLTkJAc6554JMTWi3
F8BWrYMtcGQxS+N80lAGXERa9NZezBkfr867jYoSEUd8BmY3aIiVdjDaZ2Ik21akUPxV5Qv+NmID
XKIG8/n8lRyLEiDl731dOKCRkzgZSFVuGx9vI4Q8pQ01cHUijnD+haQzt1g9gj23Qi6urmwI2j6l
JmYAmqgV6YhGuPFGcIUfT6a4OKdU7d9jKt0mXC0yjKaMeW2ZxeFHgICdGkkgA2oeAVzUwpJSngZc
BF2KMiHtHfi1lPWDv8cG75FRHlAkPG0BqiBBdbuI2thQNoPbCuhUbKJXqnwEUg3at2y8m/UXzrix
H7cqxLyReyzDc52hvfBctj6JWDPpRhOLZEfaW/gDMKvPcGB/wxptsYVFIyJqrGo5CENWaulmFFoJ
q9xPhCypt4sPFvLbxTPpQWt1OE+R3o2aXeTrr4ECA6R26+TqFg2E1i4aQuBXTNNsEo9emhs3nV9R
iOz2Js+pOHQLPH0ZbkskaMyERFa+3aAQdEJ/u07nDAyIfjYA4JHPTm8ABueglRObIc6DXqNDaFeS
aC9UB1bWEh7vqdwLwCFqTkN0XByLDL8DVhTEvsLc0iSsZmbyZeeRoUs/KAu0wKwkJxm3nCAemrC9
TcY21wEF6Y/Y1j9qjY6icGpE9PdwAxkS2IIWlhtWWl12E7QNUr8L47v83nN5PnOnqcS5HnIHwvOm
2Q3pgrllnXAdd8rKrMmPifEUYuGSjXtVydjJazPTIh2iZ+usnwbTcBfZ52rblPBvoSSYc6zDrUha
QpdqunF12JTApD/veI5XPZLjEvEN8igX3zO5j1MCGliBV4wvf2ruYX7oIYiK0nTqPhxUzIpJ00Up
9cXASZksMvY4DxIkpiHoYfffCiZ1DHjbNOLhno1kkv7ErhHkMtv9mu6eJK7nA6c/ON/fF9+hsuvy
QgJI9h3C4nEuQGDdgw8rUhO0Tc616Ziriif9K61VP9d/m27P7O2XeX1OgR6IoltOWEcdT4GV7f5V
QjkOC4C8bFXZnhPRQVYn0JhZFDto7hCslepY1X/5Tky4vZkfDlu4CQQiSTflDvIDRBXO5hECJhJO
bKZbv/msHodqN3+cGlrntiGAuXnWBGdaogeZDXKpaFb4fVvx7j6ERt1QToPVCFlYQpW/eOErQmvw
l9cKl7xn7+hF1S+H3YWDRaHklJdL+HA3yQQKE1EO8r0LUQIvay4869ZMxM9UVo8YYyy3tU1HcjS0
R+d3oyAXYDDDXaMZKclQPpgMKeA2EMsQ7yIT1AwKAGsI8/3Uv6K45BgecOV39YMthBW9cBQajzAa
ILbyiCA8KedEHUeeb73PrMEmuEpS9YcpG9x6pasBHuOUj5bD0attjZf4uN/5NTSo3SvC1QI/FX8v
dkQF0mNxfwv8I/csmUVPEfvd0iJOX9ThtzEpfS0Gvvq4ICwhHWeoXZuA6JJWAQh2myYWugdDOkhP
3ixJ4MMUEuDfqJ9x1/lvITlLSAfEi9jpgWFVUY5fZACHbjhRVlhqzryamtuTIndd69qikfSec6Or
NMTkhnIS4aBHudago13HktRrSt83VegVAR1/wcTgOgz18EJv+Wu3VME7A2a72LTXzV86eZy7rZII
iLZ5ikYfmmqIb1kZdMyc+EdEZ5O0mmy9z1Y3N5jEGcNUKs8Ki0WDR5MDzcNMJCLm+fRRQK6vPexH
HRFLdno3GqOBWMizvLULupScfTVVgvefhl4JVMy4LnZ4BObYY8FgKsl+Onj+TKvCRCBhmmKnDtgV
ojxvyQxbSs2/munlvrbowrsziKn4Q9Yv6IHI4mzin6/eu7uisLjLfPXrAmdA6wwaU03SSz8znOII
AKSjkv0uHNPuntPVJVtTzWHc4gHsG9ibTtprVbO9JwwzfgMM4jg8S+FTLpHZUT3+fDC/VpgIpz3B
aR3pB6A0X+z97rgfyR33Hlr04HxJzTadU8EWj7rx6ZE0dGItNP4Bjq42QFipbkYvkYIISlipMlE7
vpOrS5t2J8+aItljfkP+N+Ktmppo6Q2ArLMTRZKQ5wWFMRFhZhDQd6IXW/LUXdNsZzzHPflftIsD
wcaKbY9ZnwLt5zOURZXj4Qli4imupn1Kc+STXt4XjHevvlmAg1mbTLvdAnPyWxZmJxpGgVhQeVRh
3cDtAiafOWCPlL2/5YD6jSimmG2JZtMKtayOjhjti5ou6fYOKk1hWn3qwbzJDe0fMzm0Etrd7i+x
WPpjUH7frjw7DN01S6gJ/5ErMW9InwwBeOcyyl9aOj2Ha7todmyYfcLVxDZCvUtLB2vA/8w8qZ1a
QUq3+fFWmTgu9RtnM0eaWS846vslYs3GvaQWGOzCqnASGUWZscA7g/4fcZHTAuozAoSJs0UtbYGB
jfjPm+BjG3p21k9F1IqJuJMR0u8+umPHtpFvfdFty8LhgjhVc73Xl3Y/QsViCn71TZLSwPdpgO+F
eFeA+I7ztMYTVNys2NqPlilljV6JkSClXb2Yk7zYdLlCkZcjibGs+Qg7Q4W1q4WjptB7rM9TBLGU
KgddGTBWD3DTgxZP60n1J7nWnwy1ToeDHZRekJsqFSR7FoZ7G+ydeRznTMLNLrM1Rf3GM1yue8wR
m5/pnJx5j15TXE+4+31AihIKPwsA5y+3G4cDBR17P+0AkxCOodTYhc+NRxFZR82zdwnauc20Z95+
98ufXOzkxX22jsHjBiQwwEAYmg6RpIK22f9HA7q+4RPn4C5DpG9l/fDC37tAP0VBdZpWqBXIftNN
UR9Lc4DayOWmKnifqBkxCT4uuKpsjncOquhCKaxozmU50he7r7Ln09hubitPscGlHTiy31aNd9yQ
7iy8U/mZ2oI277tMIF1JulpIdYDPEy7bQq4tINUq0SYHTvE9c/fOVw/NM8dOfpYySNbtLkvYG26y
6/n7sjcMwiCNyNQNmPc6Y5OIP2Gv0YqIYPAFkB7GtPrPG0pMbtkBg8sNla8/uMDygJUk2rQ/34/x
j4eaUYsFpQ5OM7on2agaf64KQ1xDWrb3xNf4WwWovdSX1KYixUfq50jgKfjMgN26ncMpo0/YHape
hGHUfJ+Jhu11JU6x42d2WNtru+Pb+JbzCqTo/w6/fhG6/IxzG/HezentY8Xl16aQhak2eQ/LcGQ1
urIlTyja6xOa6lIAw7P2+Bc2Z5uSNw8dJQMRJTD5w/8ogXKqSjD07UZhBtL9B8Vdo+g0Kao9W2LZ
i9uklzO0WwzUouMkkCEkWInoPGm1G6nU4s3Y/s+azIP77j2JBTrXeMqYj/Miv2oqKZrR0lojEXun
AGvFbbh9Ci3RaRdNiGVhWuNR4Pu/aXmXR/wO8nv6hiIzZ2RBsIcNasMqqt42Ehx7A2/qi7VI51hF
+FFyQRtSPBBBp3WrcyBaYvanXwvv4MuYmr/Sr4aGXrkNzoj6vmGJ+5EauoZZDcjjW8LqDOSdb26m
u6tSEmbUqr1i1PQs5fixhEFHLmYGaKR2/8YJ1nDrIBjGwMzTSL8yyfJjwMlWWivCIr8NGSDpvcXA
GoUdlC93geQNQ7vJZbLJjQ35rocZ6JLQSK7/bYKTM4w9xpZ9/hCSq39uzkr/+qIL2rbOXLlNL7t1
Avoxc/45MtaqLS565J/Mr46192SEPYvWulkt4ZGL1yUvEnIAB5fYlaWzufAExkkDxHXfzZeHCH6+
VPZHAz99FQmFetvDQpUONBRDhqSp24Ff8NZD8PK2IXCPkciwz4OUxdePZVk3xPjKiIf2Pq7XGoox
rqeYRDEF0D8z/aDZw0+ucNnkJSeZBuFtglxI4mqfvHMFRrutjju29NHHGF5+BDUSbXq5WWfPDtOS
ZCKKjOkQaAmsc4xYaHMea4K4TLafOzo5TW6J4ibT1tbf8Fjgb7sg43CfrmGP9lj4J6HmqO3WK51c
tgYYD0gWgYxVcRnEQPHLOlXk2/BAx8s5rN/i0CizVMxHdG8WNpnvpZW46BpgIz/mij243Fr9eRLS
VEZjN/mmmMvavWMFwUoU8MNoW8d/jSedhQl5LHwOIBUEl8slOVFFlNlh7yZhQR/OxLn/7HSX9nCY
arqU9JNABGjm77hhj7TfBYp1BRSx1AHsX+vTKFPDF1N+5OoLBnNpkQ493Jo1vuInU+cyorNOithP
NBlyIIB+NAEb2D0f20RLPbH6pSh55LS9Lv9wf/RwBvXXjMsQllEPkdtbT6ENQQdhXcVmjPEA555k
nOD8BqU5eCxNRf4qAttSTFJ2VWJA7ADX3etyymvMzB7kdmqgnChK8y+lJMk2CfrTOYLszAwhMfQK
yqtxYOKuLMk7O7GUPE1rKnPIo8WGXi42MkEcI/hD99Fa2PUlrbzbO6gOGKHAk1BlZ4rKx29NKAcM
w/4Q1kLAukhWnsEYIQUSitNIFgreqD6CJ+k/wl8EZ0v9hpxHEaB86PJWlCV9x1EETdTkuptpd/b9
AtAU7O/XS+0J69lM9GxnkUXXjD8oXQIx5WVzKM5azmqsdnBMX64dTS9MsLyIEvS5oVRB4QsMn/OU
+Lv3tZIjjxCxArPaxsXoQMhdQtfKM+tLnm3MfitypFomBruauPfqzFOlJd+Rj5JCnRBkTYXVQAhv
bVgMyONwLgXRlpVrdz+9AlqXtN7byzIh2bWrYjn3jJzt0b34aaiAyMCDkaXxhJcI8XC/6CBWdu3G
s8LB7Bb2YvvHSOat+FB+osv+7UuaM5txa6iXogZxHC3SEiVONtkroeu2ZhpFPsHZ+YFGxDASqpnH
zlDEoNuOjoKivADKdhXHg8MfL0zaCXT6eoF2JKmzS2MksV0zvn81GFCmKPIU1OdEiPBlEOzwLLsb
tcrsOKGN4bufxwupNUS90G9zZx9yPLkz8NxWKm3wWAHARchnbgduhr1BrmcpLUDWvf+ZaJQHA7I3
mW+unzwjqlA7rf2NdDsiJEivwhYbTc1aNYKYXCGGzTE6ym9DbYJnGQQas9391Zdfnm8wFn5qp+QM
HeCEHkOQZnjwuVwSe5NXhqgR3SOcRCPbIlYBM2GxCBsLTmkgCKjJi3DLceP6xqazzU00phIIN2Pu
r1aEoGlA2KHxdGAkJQamxDcGY1LKmC+SqPAnP0xf+9qN1PfmtkbH6MGuk/gFwdTigN5V+NUt/nR4
KfxpZC41oNxoJihDpVyCS9b8UQpk3R80CRiCkDwSWE9F3d4djS2ICruWTrVonLdXKj0vwZm2bd9V
YuWmTKNmY12qgYKm7paywVPI06uA0HNAJ0UINj429gypebv2pOhNCs3KXMFrcoISesot1LDS1W/N
L0h1WE6w2gMDl4q8lqT4pZmUX9d7V8TXLJ4kM+n2pYsS83GHjpL7juGBQhNEJxliexU+1AIYM2bb
syH+bpNxUMyiS1+NVfzcNmtHOlCi6r5syCR6gHCycgrYdxGXK2tMLXBlWIUqrHwSmjSmlbRBNjBj
xOdD/P1t61u17cdBBXL5yluy9irrn4OzmzImCDd3FYG8KeHv9cbWBbegVblrchXgT0IQUMfc7ob6
oFwch0qvgWBU5oZPaXux9yeQvLD4z03HjwvsS9jebh+F+3JCR9XnSsyqzZHjwEkVrAanqWKoCy/M
wde1lHN/cuSiM4IGVT4ZiyKbQv6lvwA8KQePqhlVjb5v4YFkJodMygCnfKbaF13W1U0UQb9FN71A
woK4eUR0Ip4KjUwyRk7Bhrgp4cl6CFuQXVT9piCmPgo/I+BY4fQH22joQikAMT0Ww4bewyMGc6k+
SlrS1wk2gLvbUntzoq/u1S6McZ2iErpHs1mOAdTPK23HroS5Z3Kdx/veC5BWmnaQJkETjMxUpBcz
QjfHzyuZXCqeNXs7vuO20FI4rhhkzK+ZPxMYiVPjrEiXam0oNO6CeiDlA0YhmIwGNwkVY44MM8dR
zwgjRLCYjlgZNGWOaiJ881BdYVFFKS2U9Eqkk3g40Z+dFgYhFz/ybjdmXhXRN2CpQ+aSXfPfOh+2
j4+zdBREa+ucGylVR1GfkMfH+tb50vp34s8nXXqSdm1xyc4C0lXy//oXs0kh89pEHhx5xiDAJoqT
ONBjAiLovDuADp7/yLY0GxQp8VdA7b4gaACgJaqL5NfvZypEAuaRavkh0H0Fq9RgpsgmpFmh4S7P
ua66znUcAJLbKOzED2WzMDI4Gnig+cCpFJRMMw2fmdJQ+ucN5kyhVC8BXHo+QHR2NkYH3HTX8vW/
CjAq7cGh6jnvLWJuyTuQjYQmPNyKYtj/Vbqu90v5Psk5d621Nm0SbZQQ7Kpcrcm4suLd+UUGt+1+
wRqDQga1jKnzUmBx+I6II4bQAFQ1XnqQVt0N+pbCREH8pqA7Z5p3C+zGe304LmAmzXVPCSRpwGyi
5YXiXe47KJtkuTVE8t4CSEu1iCbTSVbJbJKUsyIbPrfCQFiuYeXGv/MRLIAmvHqxf0Czbpm5+sq2
jACh7hHqEZAQdWP7euVY1r9qsfCCIYzFmaz2BnkBYk91JUBArWEdoq3eJu/A6j/5dfIibW1gWz6c
eu17wdkU8NG+nqxPRlWBnZwfgntwUGa1t4Did+eTQh2//xpEMSQxMOzhm+latoKQh1tpg0nLFOlo
Q5KsK7GZ5gARI3Dv/JrtFQtFxKS73yw8W17wdMfRS2uNEsUsHLlW0g4fFjq+3DiG/elG+06gTKef
ZYcMqrFGBFw2P0UtT7My7r1uyyDVvtcxnzkCcijvmbAfLk/uMeQwZXyuziurxjdpKREVqyg15CaN
Jbbap2kme1i7wWC7Filh8AGus/lt146yqrDg9pjh1W4wGVIKZ5CmOithGIaINmvmNu4wojfTkDPY
YnhIcblNaglrA+ToSfIPKJAem8I6bcwesFsrxrZWTXi9RLQuhGSVr9vuetZ1FFJdhrAmx+lnwN6Q
8XP9XfXPrYytBeSTpq7p0e6v1x31XDyHwi253MrcYIGQOBIdv/IChLETPYAsogfvNggtBt2g34ZM
Z+sRP1cpgYO8rjVEQIT8R55pw8O2WKLuiWdyi1q1j3o6JrmLVUHAXDHaqyjdCb+ZcsZ2Xe4kU902
IXlBD6vTzihuzn18HFRU+FelQvhG7Rf/Ry3GQSTL/s9uE3PYltLyxtXcwQ5vsImcCRJ0metxkqcY
8J4+S46guw/TyuWhsUK8OILdfD/mWStDSwAuyswXZJa6LuoI0Q59rd4J0RLIzsfDf9qwfqCVeE/0
iTf8IeX58T0DE/EHZ2mqVkeM/36C8n+ntvFB1pQUBfQ2mi2xmroXvWUX+tTemMd+29cfKxFnTlhC
Fe0IHFwjTlLcMWZT9GBi9AZ8xw4ogRT0Z32iUR5FiqK4bPZYPONqKbTd4vm8APnGj+B3hA0diBQS
nGbdh7l2CTf6J9jA6Z59QB0OZFO+Zun/3GfxEUqdJEvhwUW64HPyjGQYtaF9eTBbplpmNFaKTtA7
1fZDC4f6PcW+SGve/croempo1Q01qvMvQw6PLWBRWlM0FHaRtPBpuU5jEOFr+Ib4lUwb4iGD5YkD
GwcPUe13PDNxdLQHvwY7tGdXbILajz5Y7XzfRKW9dIy3yQ6w9/JXh/wUXVIXUpieH9XguZVgIaGO
OJnCv4hTUXjKRR/y19v5SRDgTIkDEqb0HzxTnrCjBDBkaW42e35NR9HPhnBlDwI3PTEKi8eg4Fpf
jTwBglxsn5zObITzsN3HueN4+k3VQ6Y8RE9GGkAvCu1+Okr2xV/4EfhXz8ZRU3myhtrimzy3rNRi
DZxe448lCSXT30TEDEk9LCHqSR+35APKhRFK854fujC342oxhFO39ZCf2DjOy/dc7bwnTp+Yaoe9
LwRnLAsa+q07Yfw3i/ncDkS/VcuthvemxZLcsIhmdPAYrqngKmI4qAHVxMaVAx+uNCP+6GPh9XNM
zzvpPgfuHi+0yTlLJZFv9qoB+WCJQ7ZTTGXuYxHieMoGqH2MwLFDq1EBizVpZDgPuO0vNtvFDJX/
D7wiNj0OUY1S/y9JmtK1zirgkt6gz2FhFpxetUMjXhmRkhMpmxpIOWJWQZjJT/DmrvGhxSG2d8Dw
L85R5tCbFQtt5SNbGHvLizEMjXt2Jgix6CVtuZN/irt16GAphIM34MujmI8xA2nP+tUdE8tS9T1l
nfUBQ6Y7g3K33ovUxFMmTVLGD186yuh3mtZM/0B9wbCuUhW0avrNwYtXFiYc0Q4nimi4braJOV7x
9iYCLgIgUWxUK82UMQWsJXmGrowgngEwqsCJd6+jjF4+d3JbcF3LjU/4UyrKO4/vgBdKSkKvDnzn
PjjWUXlCVdMfdapy9wsD/QfvecNqX40DPvPYDmuTggxXPJlM+3tZuUH4UT9rQy8mie42JbNMsVEK
Y/x1EMQx5l+m0pBkUjSkdJz1TqDrUThqbiAqgorkgic+9xJEPXKQQicuUbAx29IwfUYx3az0Qb+4
vvHhAt7dbVUwvj7Xva3T03JywLP2pBKpIUXMavABXTr5SwkVrxdyR4KrMVmxCcGzt+lI2Tv9kP3e
CdGv2v+vswxqobOoLVQsHfoEUV9aIXoQn2k2ppE41Gp9ibwqS4L20+4eUiEyRohF4K//fn2R2PNS
O/YBIXU9Ep+m1Lo2QMZrCNeyz3tdQIp+5dP/DSdOga+uSQaOcauYSa3SWdUf1JAVlbbPfDxIP7aF
vUdNb+uCqUuu+6yAJM+iL5zk58zcf2iPoaszCfuE4toBxzZAdC62ElETS8KnHHpKnlbh1Ckijg4R
3DSTkjB6yKpDzF0GHhMDa2NgzvwDvcALl03RyVlplG1P150/MAjyDsALGiOUtGWWkN4nTBQldUlQ
WtKPvVpf4olqbjP6U1TOM1/7yDJyGIbGDXtdOS6XZmgPT38uvtXSbLqexGxVbHgUWgZkRdfrj61w
qLZzrTjvQGYhZMvxGVaJnYvss3H6+rcrAlZKKlRX2cEoLzRlmRiWYCnuvYi7pPBofnkRqLY6s2Fy
MxWP0FDFrm574oK9ncgzeXOUNTfGra+/BGy9nIdN5nNiH2u6Q7s9/9suqKKadfkAwiU2ba1szS3K
fNvZMTg6YNorGSzFZycptkq+q8CWhsoDHWOxV7z7uQ7vWvOJpD1gvaByppTtMxSR8wKAKtqRHNjS
8Pt4+Oeu77gDXGybABId2zndrWjxqlyDQPTOGY2qr66dPaW28Z9Q2ijkU/MJOR+rD33KyvaE5fNW
pdd5+hDbqQ3wO/KLQjOMU815Xx2qQXrYJpmZdiO7VTmOifduG+TZY0h1t9JDDebyjYQgNyVuxJVB
OwIb5fKAYqJFsXElOa6OytEbPZvAPZ/M9G2hZcMn98jJ2qYrOSpNgz2+poolIvO4TVGE+IMxL1mS
JcqhVt/zVbPZCpLmq7czM7rXmGM1mGCYS0u3qgGEzYJCYv2vZR2wJUcnvJY7tefHCMyGs9Wo/ols
u+ALCOiRoneyvwREdrFdfLUjzIkDe6PUc4KuNn05gRhPCpMjydRTR+bLSYXVEKeEQeOUQCIXVkbg
2D5oWnDk4Xyy2gVYb7JHeOQDvFWTkFDD9ZZkNlfG8N6ZEzhJn44o172UvmNgvwCv18yNEqvlD97A
oiOQMBXBbCuBvBXvZm8rAI+Jw/qfU6y6luF+1o4baUHeUOd+JXCCxyNrdLjaood1KAUwtcUHBxWg
AiB4vnxR6XrAzbq33glktfiIu6g+yl6rCPt+HF9H9S1wMngynA4wJH5NsluH4/zn6nsLq60mYMyu
oVOvtt54iYl6drNpdNTyI/+H59lcZnMuaAq8v7ZHI92gwheVAkxzUespbfo8dY4NOQEQhgEPV3CT
37bvIx8oPmKOkkgoIhPPonusSEX5PM1mD7dRBsj67hjKjBfGN0glwxqW8eZXe0ArYCcMU9t5vmmt
tNxg1C1jC3JZCjbyKhBVE3kdDHB3FIuK3e7GHHmIa2wCECxkbAZyrZ029N+Vs2rTwP1wkUnOoHvO
O/7nTOyHhOspCQGmMof9mMV/vP/ko04sZF+cg4cdajUKsMrWlBFyqVZsipsy9zHfHHsvI7Ehd9dN
6uvRHI77GEXmdMag9IeI4PNZNVUR7yH/3/vKxm/11Ajwf1zcC2UYLDywBOpXYNVPjk/Mse8TEFmB
ie/EDcB/uIeyCj3KlfqdFu3A5xjiVp2qwPkBhFAWckk17mteajPCyHz3DkcbSUjV9Goew/QPEd5z
71Yue0YBZnaKBNkqspWVtDzPcoykuCVxjhT+5ZNKgZc2ZW55vae/UyybgcCJSvsWDTsqc2iSjdRn
JeO0s3ytvdzbI+2DQL1znlmXPkTDnvbW9WvkdgCLwEUHM0yOALeUtAgZidmhA/E+yNJ+ev8+Jk71
0rS1MuYC+HfO9/DE9htoai2TyjPpD7w216CqxSAZ3m9LY8wUrI7FtOC+vrmgtGrmRiZfj67rzE20
eSeJ0jif2JE+YVMqwHiwNwsH4JaySt3bm4lrWu8Cq2CsQA1JrIrTURQDcdwlkNlq+LSM1D4JrALr
ABAKVIGqjLp5K+ORSR8xTtxgf7OoVl1gXAsFav8xS2NZPCzk7GqmOPMd8ipSf7YPl6zevWbTqaMB
TYBqDiS92GiI4nNG7EqtS/c8bRCmvQvqSpumI5jFtL1a/KflzN3+z2K5bByJkEtJ0aHN5BaD8z5o
+EHYI6oZ32GTQbMryYu7eDxG17gGQXtOpn1ZyH+HKAc8+Qqj8uN4XyJTa5q2+mtKLaOwjjCc+8Ok
vnbxpP93uHOKyq2AY59nFMakhixAj9iDzTCUlGvz0quN1HXfmUZtLhgAvYw/A1GxZn6papmikn6e
mcaEYKTjJWzC7yCP6r7Ym1wK3bb5b44BlCNdt4SPncPT6/2XjR3DXCu/FIu61j9NUgrCwIlovwYF
AhIk5yPd0wbW3HGCheliGP01cG4kDVH644lZxkVh2FzDej0mT9+doohka21Kr8tGB5YaSsiykaAv
JIQqFvV/eanKqkCgEoBqPE0FH0/Nmj16xnNckFADsJwoC/h8U1qOeHIqtnKXN1lgalzov+p7XItL
WYRstHbjMtlPME6pGykIpKEfmU+vQxYRC8Imn6+PuIxhaGc8arN1ch8o3e6wOCdAvY08A4tdOIqU
hQmLgD8w4chb9mef5GeOlUVopBKneMtopBL5u3ceSVUOh9NtrA48jOCN79maoQhxsvtnpfj6VaFu
zgadziwl2VQTCYd5WnDfamT0/5t7crBpHE8DU97Ng3jHFLlLQgKCGh6XzvO4x8v3jkzhv/tICt3x
KmLEnt7Kg8lYtCb0QIE1OCEqTGCGIuZNuHo11l7fKjujaOJL4aq78hPDIt1S2sIPH68n1qQjhyxN
v2rz3cdzukHvnIFVt6lsDAz5DxHQDTsqsTt1jNFf95dmOFXt0PmbqaNFj0K9U3ZoShaXeJXheIa3
i5nK7WPGFEIE25sLdaAJ6fOR1zGodeZsOMq0GhSLbdbE/6oCFfaW/Qv5B/mN0EY8HLj0Dk/TqyNz
yK/HPcvsdy9nCnUdBBknPN/jNeoc5iR2cQpZag+7zdcz1hxT/KH5xaYmw5FH5UTf1oTNb0NF7iq2
W+JwPssEK1RKFquLaboqDK66bkcJhdkU7XvrCv4NorXOZg4Tg2rmF/zsLZ/RoSV9IDZ8pgsFSK/l
vcG53Hh4Bz27+FvUPmPvOb09xVIFPGfd5K+5G7qA0v+yNzYTNkSUqHwkTRGxChkVWwvfIXRXVwWr
2a57QwHWmnShjCqBORwARtHabB7kcUJwyYdgKey1ovRy/u/Dg0yfikagUXaVhy/XIoCuXyBxzSfB
XEjdXS8rD+ryqG7WX7+Dn4EeXzA7glum2BtU+9KSdhgpICP6zGfGELCvJZLtcyaNj/65NizQjgWl
ikmWI423EqUMkeGRKgKVzart6Cqajxu6938gY6RsFv+lZwPcdg1YGClBSGCoM2pF7E1/DUKGMOqf
e2uDbErmyfeNE0BOm5BXXOKr968oPCKQFE8x//YKbGXgTXEkdJJLLlsGAhPsXSwX9sLRZyVj+9He
lbj1uFyEeQlF/mMx6tMAgcnDQJlhOxuRSRNYGeX/3RJPahT2nDVw32HpwHvwf2ZDkpFgUXmhFC9J
0KEVOFbDshCrqXD2gGNFWsAhh4rC5Gj/OvuSS41BhA5gNvgHj65LSdCeljdUAxn7bWxD34PSefjH
i8sDJ4F5+J6vU0UD+Tl54N8egxOv79SpeQFTPSDed4+FprPo8g3n972kZ7X1DadP9IRl+g67gwnf
5/AvVHWUik7qI+we5j3FeDJdFzgJ9sE+LaDZS3Ox8cQ7olzgpBRLWG1/FkQcPfA6mjuc5OiYbTz1
4CU+V4dPYCc5tWILdF8CHnlIytSlA26BLT+8D9Y4Mxc+9HIq4siscqXWVh5pVWQ0YUefTl+lbAPb
Syx6RgA27ryfH3hjBnKlh43C60828sPVjDGsDYFUj1HgqEx3ItTkiiFMLZD+H5IGXv6jB3Alvxx7
mZ8lrihyPSRbIaRflfNyO5qI30qVqxE4AMipN2JRf2RSHgd9UyYCnFZwUhXgmjiPFb9AQ7do6JUh
mb75A5XzMenDecZ1Z/sCCTK7lOrX+KR5qK/eq0eBXGSSQU7hNnpxiIA8mbYL8O/axPXqXp726MX5
iGiTRkphWamdUJcmCbKeH4Dxj5MwKHhcfJNDU6vBdCnxkN84OmUkF89BpION4XNGoVtok+1U98Sj
WSL4hO6c0geAYcObJy+4VMedl7XIm5qyiVXy7nFhYHmyzs1iJwwNBZ5xgcG03UmYK+7eB0AjmJjk
xkrkcdG7kevHHiMflrI+eoon6CNSGQxHDsQqJ0MUHDqjNo8j5mP3JEjsKiczS6llAsp8RG7zZqZr
0u0DlfscOyM2haGG8ngn5zGRq1128qLi+zVBQcwlfFMA9lLHxkxsanY/unizl+pOvJwWF/JdDLKV
FTg1mLcJ0uYFOadMLBwyL6+nK0UFZHh27RG3TkGvxiZB4E7p+kQHExBDV5/G1j3bG07zQILiQAoe
q5jqu1x+n7v8xwy7PlbnOK/UGlL3+7RS91jK+cDXNqjwg6gfgLg5RbxKzbs+YIbaaftihFNY/8Uv
fA4pzRBEz/DqfTTpOAhsytO70MYV8vTJ4GgxTFFQ1wiY2vXVeymom/iAohnkEUX+38l6BoMC44FC
RcBCYALnow28Q35usEZRtPoepx9HQM6XN0gUdDUlmTMPkToQJStI+Hv9I/M6pncvn9/5su79plOs
xna97Vbx60oEZkI9ZfRxnW3s18xBLsYI9nDOqhPrm4RLLd/d/AJ8RcsAm+NrtwR7TzcXomAgwr0z
VWHZ30f1/b0ANt6GDcsZ8qJbgO5AvwkMerxKueqN1jdwIhtP9YzK/o1K8GjYU3IkLAhm0FtR5QzP
TuYwV14AqbVbcpZasT0Z+YTQEpOYkoo0I+2LI+U5LPjOdFaxh6Hvpn07bQiNhWdX0Cyg35pIEJfV
jAbSS1aQjVDJ71hG46NgxNeLDlpH5ZcIWAYqJDVwAdWMwo6fM3M9MGTovspePVG0jmt8gL7WSXSx
/9X09VRedI5WV26BAlZf44AysoSmKJESYBq/Kbux+Wz3JdyO99elQVH3qN4C089sVteCXZpesD/Y
Yt8bUA2eQD/5T7CcEmpWFQlDlhybsS58R0DWJNHRqnDcUXsL+8/ab+l/gjMGu0Ss2O/GXtjNXMI+
K+pc7tqn7aOMsM9T5ZyQf6Beb2Cx5wGSrszCfhnRwKgNfb5Kwkf+hsBq0chF/AMKer3zVTaLoFmA
Y1T/smISfhGu3lgWW0dqRSOxHEYAFnm7sb1rtuoaDuDS2im9ntVLWq5PzGCdOBeAFCZynVS7NTcm
mcdzYnHvv3dMwxuXW/Bah9QYkiwzYh2O5O9ckkN/b6QQMbHm2LehejxhxJCJEiQJr96s9C1JxTiz
myQjHIeY8mDV1UISvLoe259yG75dC7Dm39CfmkkSYtHrLo9yzqzYWLLO+M1j5rJ2+D2zi5goR+YQ
9hvoH+nF09ZhIvEtZndr7ZnsP/8V1RtXHuuIlplVSEwjmBuZWMD3j+WnKxcZTUQrSpZi2wF9D5/m
zryJ6GdBhCs014jot6gLMfeSUslXpTl+jcijXD1PhelPrC/RNS6KWYei/cjE6ao6sJS996G1hFJG
ov1BBIpgcg5xZPmTYqdkXX/KY6Fvs3d8mnnMBQYH7xCxV7lz9/ZGI4exTs9hutjtocJ4QEHOeVmQ
7edJLgClpPCUFW+IromI/Va4R1jTFgMrUJ+qEeCRXRpCmGvw76St5qHVUoQYaJKB++L/xppABh2M
Hdsu3zRkCeHzN5oY/GQPS2NtcLZy9RyjJ3xALa2ypZ1/UV8OGMQAcNsIcNjFxujc4gOBuiOFj+kX
0PzYB9uzIumoABcB1toNS7eKU7bFkXPxI0hlD6RMNM5BIN5klp71G+GK63M7zJ2Znk5I6N3NsjX2
980sFrGrL0kHvp2FyU4SSHAskyTx9dzAkEF5pMCJoM8EMtQQDd56Iv0BRNHh9fRBkUWyvq7T1Siu
CD1abbrFTfx0lSefq+bTLZ4pEMo5T6hWYEY7MNYNmRtvBx/Hch7TSq7Axj9y+v2s0pAUmcySlZm4
kLxO84+Vgf8DUt7AKQvbKutvUEtJWjP6MEH8dURz1LUh1R6bN/2zEp9LLTlDzAt/6QAHQrtoeBTP
jiS3eZTyQ2vSZ24Fwr8oNQyOpiTM+VnchZOO1143zcAE7YfBOVPDI/c8tui7kyU/h6ENpowwWMCb
YkD8BoOD+/uT9hYMQv4tgZa22iPLkbkoSN9yhDcaxJjr8CiDhlx5Kr2dVOG7gjGyWHcvI/4d5/f7
7ZMBo00l66cySuT2mgaEnJsk4yorDy3G3fZJZJNmfKqJu0zqjYQOgRwUNaKgL5IB/4mikqS/z87G
WatY/iGE8DB5baPl6dI2Tt27QMvdbA2vdot0N3mHr05D2c4gXnv23Zl8Ra6Lg6LXuXwEVp4/mUD3
KvOEORO/tQcRztnzIdopjEuYFLJmcKacVltO5/nLWFxiRRKgoCdOsVEcAxdC9LkcJ+mbqOo3eCA0
1GSmN7xesPfnkRj4dlQlREib1PAT+b6Q2CrGm3FZ8aT8zSP/cH65fmi966UEMuvLKFVsyp8h1X2B
Ax9Q/s5bqqazkBZkG6NjJwa8k9YDOYO+80KBpFk2XU+mq+F2q6hAo0M9AkvwppevUwI1Chp+kOB9
o3aUVjT+i2Fo/c6uiJqmxHmqLC05ASuKOJQThkSB241zMl6JSp9yT+5uCrbHw+MX2DhF1YyfKssz
32noTJDdq9JWizih6Oo0NLLqX/i9KbS+95pfw3c9l2ZA8sKfsy6U1eEmOTldzoGuoRvdgh10MshE
6EaEXcFNIkKJJ+8Ha1bCMssPUjSw0U0HkE+TdkO6z1SJ7SotsmHYca1WrH5GO/hvH66uWh15eK2X
XPfKBJqZAx+V40RjSwqoGsqi6Id5NJcG1jomeQ+iL1/jTRnZds9eROgq0IB0DY9rI/V6uAkKV0PA
1akl0lbXTs6gJTzZxJ0SGm6gg4I7orYJ9h/hBeQ5iBAsz2y3p15kG/h82ww3Dr6nnTUM9A2CJleD
jRMpCG7XRoWaDxZr3eCgDjWpKdW5beY+Ljf2GnVZ2pGSdXbIRhk/E0zF0xDPtrkm8WG39pOChMg2
YTupLfJbkLJ7ojQQXerAUXWZ0RNpR3YJ6aynSW0YOFAGzjhygsxvRPTN3C8GIMyy+Ki1BbPYbhBG
fpG+5TjNGthNtuud//FsyqiwhjnuQLS9oH4pcEI3sgqRxpPXSeHXhsYOoO//UrX+d1VfE4EQ7z85
jTR6nEloKUUDxVY2FOeWM9UyOJNZiGh3EteUWupIhRGVvdKMY+OTalzrJ/pQ94dVTNC+dNP4jljz
d+06bcoyfRENhrVijfaPI6kAmBfTimFrsBj7zgoFVeg4cmovYAtBR3NbXehGExvTCESjiu3EGBjh
oLLi1kod7GYX5pV8z6Ej2nG0wdzJNE8CoUZ2ZJ+3xV9x5ma/SbcpqjqnBK11Ehp++JC7Cz4ffKTE
PBIVjG7XTEj2BsMtOalJnb6AEFIc/+ribQ/aTrTQeMnRkSdA6svFy/Q+BPHZXTlZh1Z2Cip/f6xA
TLMJsUARF5r8yugb/RqO6tK6wLJX78LzjKE9XNOWS3OOTWDzAl2+k10P9pLT8CYDci4dvYjqAgY3
J7ikC71PPnyiPOfO2xstZ8R4wnwuu1Oj3MtXrYp+qh29tNmhCytX7D7Z+nkAm2+9fPgI8RffN4P1
mnNh1v/MHDCHUvFa3iqmjdBwLV0/+Olnos8J5lBq56ecOXbexI7OxtH1Vha20x1cN/eWegYoTORx
yHmTCM7FAChe6OsEgV2yqSl192GnhtWWpYGn0xymag9/6fHuKvJxDjQkYPVXE4/jASTyeHanjq69
dq4EisA02sxTbJEDhylGSBvvsxKCOUy0fxgBlX3ZIlQcmx0CNIowVrQgNG2XGqeH0Uw9A1WrFDqZ
pmBP1fpeJ8qjiIwBCCg9YPAKowc1RfepJ/mzoOeTfSkoBjv/2bIyHc+Dbhgoz4I3Xge9S9iynCI8
72tKi1vdk8Go3/IJZPvcrMD/vYzVsGyjCcgtROv1aRrEBOsesGNWg1yypj3kcD5vM8ff0JzIC+3X
gQgc9nITiBImYkomP3JE1VJBq2s3ouQU+irpPgikvA3vHozr+LiKyEWJ5D4pLUDkBDQLSxOG0i7u
4yL8LdpfVk4dd6K+BjlBJrImTqGuWNCG5nJkh9ATGjY7HDgX58KHjm2auWd9YJZCAm53W1T43TBp
W9G/fAA27mO9AMLQDMCvfu/g3rEo1b8VwA5/Bb/hqkVLifMk4qbDxLVJnrTzv5Lstpsg71sCp0Z0
nJshwsNg8VUKwLS5leV0uJqtXWITP/7u3cndA7HvDGkGF9SiPRZwGgWUkplLLREDruBuqp30BLKR
q3nYTwdL+3D2qBFPBmJL+vkMpbK/ZAWdVVfMCgtQ01swU+0s44ba9KnGxWoUzUV1s6ShrnSqlGyT
myKoODb+oXl3KVxU9Tnv+Vg2hSs4+zQwaPQFGY+Z9Af6Nq8v2+6KcV8aw0ecZLcrU8S9veJ06FRn
BhUMxzMqi8lw6LEFo/WmOAxXeGbe7GHMvFfatWoKSeRjxLR8d89uTydjB147dfU88rC4bNeVk3p5
em+T3S9u3QeqAM1HVeaztQtR1qqdnTbijOgFjFN6Pg4KtO6TyfNfJ5KyFv1tXVM/VzP0rsql1AJJ
mcKgnGyoz+FstM0CkveE/3pwXA6XXo5qE7dpXBANmo1w88SaXT0olWMOjYe4mh+eLpPUWGB8nr8/
qzrbHvgbvnB5tZwisFIyK2HzPThtvLTuoejUvZMb0oTrHJNn+UROb8+fgqFMQcmnRoGBZQgtlj4b
qtXOQ49oU2i5GaKuxo5YALe5XDh7h52i0B8uq3A0QfHp9pug/X0dkeuv6Bb3aIXKkGrM15oNdx3g
cpqIGwtr3UdCpWlISOqjEMCSykBkVSvxqQR+vk8fPecgXnNubxJsQfY1nl8uDJZXxnlB0nYrHljt
SbHJr8o5EE8EFaeT7PxwTjATN/tw13IDv+bU66lEr5U2jntr+KckMtvTUzdqLGBmZ3BhWA/7S2km
2WQ9WVvoqvuvms9tzAsmR5u/90FybY13mFNFvO7ezaa5MmJ8WGt7rpZmEm6x2l4twsnhLSZ+v5ji
wNlsnoOSggbwCBE6rNdrkIa6uyoGkoe2XtULpqDXJlGtSghDMbjA+M0SN1Pnu7SqnrRhAgj/dTkT
UcLc5Xnh2Xb9Bcc6GWoiOAYcWaURhwNi+sj0A4mOf1SfEkDTiBj14HnN89NiQ6w5ycZh99KUvzQF
NTQXespwM+uhLoZ/o2YKkHeS9e2YLaLz26u8pBVSSB3cfUKboV/Eg3D9PL9WTmOhUd/QKKvLRLCP
7k35qGu6OQf54Xme2pdXKzBnYsfjErIOog6BeFoVgZBsxO4s2yFt3WDOBkjSG0khqT2lF1KaljXQ
l9/vi0luKwldXwWVIm2sirrs06rCUvz+QO/j3+dF2UZMCCqauA4FM7+QKG+ue8lFq3YygjrOCFYl
zLa0QZf+YjtFaK0cgmllqya63BHEkAILOZBB09ELjiwMwTfm+ZaBDfVNbHueiJemds/ji0KONIH3
IJNC4fEl/nXMlOYxmqp2pFt2JZ+zP0AjKJMwy88cAoXp2QVA4UPHDOEgZwnx0+oYW1SYbxoEg7HD
QvNxTOFjPQj4WjHEd/9xLLPTre8WXDjuPbNkpsxX7RCIe8krK2u+Ke9/TQum3K+WyVixHjhSuPJP
ZPW5jYzePne36v7DfVEyH153qkCyjCchTXGlwR6ONgCtVeiOnMEfr8rIEh7zzczy8la5NxLpiyRQ
NI0a/Of2YKXxj+aP0ZYeCzuHeQBeT7ul9V0/jDMKIiZa8PdOCj0sx9rtazc89DRnbe4P3CnA0b73
rn80NtvfeQ6nYNyi0H3ushhW70EAdH5pfvGeu4tb/NW05vyiOMh9SMCIJzPA4XhRcoOTID2cdiHl
wic5krf0llKR4AEU9P4Veg80L846lmFbb94VMYhqwgfGT0nT584LXOTlkD6eXpsbf2WFdjhitFwE
eoFXNx0CZJD6MVpaC+ttNcvC4rLMaHrjSal9Wogcud/R5dQ7mxk2dlHoPYgh1cuWk4XV75jFB5QV
/BCsxRETBIn8BrOuzDoj+u6SSiLAiSfiHx4l7SLPPzJ0nG9vWBHUpE+Ng8oW1rz+ftI9Scqd0D89
fiqq+4mX5qPP0a0dT98ysN9e23kfMc/Is+7JCd7FuzJDlBcnxunS4Z16aiMZ18QkfIqR8i4DlnYx
9MJovSXSKBFDVroaeY5lsJmSAow5twxnEi7XophDyGBaVtkx1aoNo09+FZaAu6J3aBY7ZPdegswl
Qs/7dTWJ63RmkW4UR28NI/6n2ySNblXpu/ovyOhaxi7rG9nEdtrvEaNGJ5AlqOovYCd2TR9BDJO5
tDDC5BX82K9Af9uKi1GZ56NaAiOkUeLaF3e+mNi6m9ASYTmwBiO8wh9QtyLp6Fwv2jEYgHA84Qi2
IygD6IUG9NSJzuLUoq+eebO9wl1urZGWSYDlhoFGgd/HfwFBW9kYmGxb2DryqK+Lx8uBGu+eugUz
Gp8+qSbDy0jHBgJSQxVl0dLEfW/FHTfY7jKw8odmmALynTQ6LvFsN3SJQQEvfGBgk4dZs8mD8GLW
AuF66MAAYu4nFC/VHsSyR5KM2bePgh8lgSLr3pjriuaieRTyhNdkkCAtaycOse4JhaBLwe4MnPNB
kYsQLZ1WznE3DJdtXZGIRq27ahhEBOqa9cATG4N6z60sxHFFxANrKTLl2e/T5C5LoBgTkiJW/iaH
G2RUXF37tdIm1aWpsfIyu61bbMSoOeuC36iOoFaHq7/3C4y0L95CQhtmxVkZVFXdBhUGJSuMHDdB
+qvs426Rxr+sfWRmNe29jkQS8xq6OHtChR8Y2ebSaUJnENlQzbL6enL1TRtXHDj3QL6/A8YsgJaJ
QjghHyNHu4/6Ik9iZXoxxOUTDZ3W1WpJMu189spcLhevD+MHhDHGqrCPItndjN5lwaSTpk2Yojza
LLfQp260a7MuJlPy8UMgxpOk5W0JMgiEBgjacVBpqBY7MkhYQ/Kw0cQRYo3j4W9YI7ojKdruEapt
eUhhcwt5sBospgTXFQ6H1L1SS8GXufbgzNw05VSB1p9T4KChTithNgmye41sxSGhDb/Ezr3zWsYF
S65ZT5lAmjjt6g/NmPbOF+Tb6aCOYBiHDnrmpVUnHDMfBSWd49VgIgpnrlZGiJQhHIkAUXuu+s0f
HA2GJd56bd/zn+hIk48AcRWEFvWkHWAofc/l4+iFcO5qd7/t+X2wi8QlwRD6TLtEUSY0YAF1XI+H
mG2cENcVkmL15iFJqaZ4NpP6LfJYmH+oHOMjZHUKWRwTxmLP7W+7UOeMEWk8YzP4HMN0alkInPAJ
vK1GikCjGcWOjthq6R2XBzhiYPHZOKot46FmxQ0d+Nzs79epDDVamscIeEjzJtKrCGGYICgS3/fU
FF6xivyGUD/PqZz4n+i2LMIbihVH9RyISEJYOArb0ja6opmDQV6ZUxryXmgG03iw0YlukjjtkArM
nTeN/IaDXq63OFkRqqxoqR1tVxaes0GPyDQ3dM6VYaUzwJe3kWZ/q+5lExooCrxMQ2L7vxB2i2gB
V1hlNyRtWVoyDA0b/mkrNNCRBS0tNqV4Utu4knt9UVWQLJvvYgeDSQwI6IqrRKqWoMRymiCKmjI/
jDrWZEU/jHpa6dDRNBuNKhcPvX/uInSduIEdP8rzWi5p0w9XrfpOwpVl8KJN3fuD9H1OUYLDEc/1
lwWMIyex2AUiZpW701kmsn51zQbmTxrobW6QsTfkxHF0qfCDsKAIzQWlBfkuYn8WKD0SkJ7gWmx2
t+pvCGawyveTwxPJy0xSA2BqScUkWq6hIWV9vrQ3xXO1VphI0h0Ds3Hx1vxt62uKuRRnXS6siRZr
7lAqp6lkBz0D2eC1y+g2yU+KIZfSx/22Ye1giyzppjS6j9Fd4i+TEIOiTIHd6tjgKviFb5hqhs4R
GMy6u2azo+Lp+D4Y6oKhXyqH+lzQDiJjfgq88yLWGJjBRMWfEu5ksakCMQdCxzL9nPYMez3tTY/x
VEi9ipKfxKulAJnJkOGXE97T8ENhH+z8tG5bzMzLyeVtpGwxb7RrAGJH/yx5VrB57J/qvBeQLwnl
g1tHaYGNI1uiZovoQ6w1Hofx/KY0V7wxHBKK4hgPyt3Ltu1GJwh5Fg5sHvdcplbI8SbrzR8v0iPF
6kCqvPSQqx6wHmoASpXJpvNgqAHwD9NIhfwN1zWx3bj4l8oLDmia5F1TbDMP6iIfu0HkoDZ0IdCd
1L+yRGoeIlRxc/52SMjQc0+j1fHUPfG2+bzWM3U63A/1+n3Kg3wZ0T8UONaUsdllxTF/co7ARhl7
AtHMCzgGstbfvXZHCZlo3GdrcmhP9xkMoMBS9O70DMDalX77E7OvoNwYLIIHKCvLtjUoOlnTigUX
5usmtnceEPkA1en/ZSgZ8T9WspoU1Cz5QCudEwKqgRSGsenl7JfxTTblpVh0hYJCw65bYH5tu2OV
UXJSR80ur6Jahf+UP/kVbRDTz/dSu1B9bZp2S3Hiyq2rs+uRGTT+2ZEt6atkwAu+Hlm5gJw+MVtt
WtCASNLw2E8osf7ntSaPhQysCpSAHutU7hfJ0N4jsS+NEHmsqp2Go0zE+b/Zm8cr6Hu7+YmvDts/
dDAi16PTrJIaFlThiPodRvsM8i0rl8y9+e7wLS+PUgMKK7ETEm6OgAV16V715j2IkkituW18VWVz
Xia/hqB/ULVtFy47w+lk0af2hldp42wf/u9kdTV7r+bW9rHl/s4Qfx9o0MHRMWTljHW4UeKU9gjT
0mvmsdoyaw7yL1jUmw8c160t4bBz8BocddzShE2cpOE2mIrl7TZ4pmXvd8xhYxgoasclLE66iI76
XrqWPyobkmGAx52hW46dKTdG5JsqdNtpGRoT3EHZJ6/EYjcykoLyFDKzS9pS/8tMOy97FNl57e2L
56JPb33//Conepdweb05oLtyE8Cokl75af1wNz7mdjqKDwTIpMIgD/gLyYOV6XylIuUSpRDrVNpT
Tt9IJ7L3Uw/jX778X8n/hoe3pEhC0CKFbOiCTc1qBjIcWM54zbnV2saS9qSJa6BjFJmbZIbe+Fms
vATKPhkO0b8Dq5qL6WS8GjYqZBKSglEpmaQmVK9UxKx72qolKQmwI8iTi1br2cTOr22ZkFDxfMXc
3+rSxxD827IsaEEGxM3nx7vwjeO8A4mVZKX+KdxHWjqU4QQVbYsDED2mXLSQW2kJ+FlKz5RVL5Tj
SzMucH6KS0Z3qJVgd0oxNxiMYhxBZyjLqZe9oHtVN/3nkEG1l6y20nJZ79WfXLAgO0gFALDK86H0
j8pkqR3U3Ls6WAfzy2GidGIW9u7YTy/X0F1k38kJ0y1V++6Frxqu4vL3PuSS4WJnRgrygX80gcHO
iVMxeUKR5x3lQSpqUVPu3B9o2HUz5Nr4ziQ/klUT+FtkFjZsBTOHijLmmOQhXPv34puUZhA1diUo
qplmsaUKsKJQUApvRdkDrRxQhYXGOPAJ/efjoly5NYmpBcQQPMNLwefvFr1umC2Pn2Q1gi3bIwAz
y1vn5y+c3WNOwQcG3zSF/jVMyWBfYsX+0Ao91M+65Ka1IyUuQO68X2GzQ1QKaflVzzGiYW3lOz4p
XZ7D6BY9EEyRU2SoinCwyp3WR0XMrkybrA2gDBhWFN9bN+teITZYrJrNrasLG6XEtKIUm9J5hiy5
jxRrV/zLRmh2Nh0HQnF50i9NJRlIVGW2Wxf3tmN9GyGl4il4HjitinxiTfs96wmkRCeE4aatwrja
uWArhUEYZhw8fiNnhBmuhVbBQd0hepVvH3f5w6ROqsUcn0o+j+9Ud4XH/FXZEVLJp4RgabwJLOxS
MUx/63I9evauMCXwOo8+lWWE5Ohro5IczOJBkpGY+8Bd+J+ON1lMVW+fKeXvJLUVrbrewAMEtVC0
COoo0rf2TG5Bz1bwW+miu9daLReZueSr5MYWkAqJH3GCJUbKlFOHYya0CGuLPA5MhRy824hM0Eh3
7yPgwHrMLP85SGKGS4debh2n8yjdj6eN9ijEzjLTmQ0NaLdNtGyU/MYmvcYTzxkWqxS+0ZOq94xU
3+0KGBt7IOAUTC8drnKHfLxOnfKMGc7hmgEltybJkhWXQt2uaPeVjal9qXpezPsT1ByrXzIm7gIa
wHdP14DXkNJQHX22u+rM14PLVKz6JPOqji2VMgPWG9dZPT7bnfpwfFtqnhVIfNCD7tKWBFaj8wUu
n5Rwk06z39Zu7XqCH9clq05QxU2ZaJNySahCmaIABBqN45vHBMbb7obFvbW8rgfzyMN9wSpQEfjA
zgovEJPdKd6ElOns51cMyc2n/di5Dkeo/02eTE8j0qIsQ2W3kuXjFS4JqxEAu0kJk/nz14lFmTmY
D1OSiCfQOvyCbfiLK83wvF6AEh2QxRV8uAQWGkORCtciHRMPhmEwQU8xX//EWKfzL9L4zYbXonGS
yxEGT+0UOmPC2B2NePWBsVt7Mb2wgiEna1xX7oJzYVmopM5CQRrFP19XyfBHINRH6xrm0h7VEFsR
B2avE1SYAJyO7QU5WGLsLEgvl4vP/wjB0drF8F4xpYK3NV6JAGjey7GUuvOoaqUdk9TwCLgHedY7
G3XJdsrgHDhkpE770LZo5GlfAqly6ML4pLsGflN5MsJNJLL2iY86A/U1QIf6Ew09oyphyur4xecz
yoDYTW4Jwvf+kOwMuyFKN0D6Xryq3dnY/aehjUDAMkbHstCPc804deWsdfzi7BRL2iGpZpYcsUXx
NE97HGeGWKNyl8HawUAvwKUr9DOZeS0rIMcHEljtxKn5YGJyb+vNVYJuWBCCHm54Ek4hIhQcPjV6
VhJiC2s8RG9xtBxFWDVqzsTbW5tk/nFx2dmFtlruMVGeY6Abf7oNUakHBIaPrWB3MXDX5k0zNwXi
de2gO6ZT3ShvuEJsOEFF7ysZYHAXn2k8SXaH8HXyFktWTva/P9ztlKcJBbzwllLJd3RIVILIbRzd
EdZPnV93qSwgQXczV8FbhfxbC6uAbxE9TPl+QvpHKLVJMbsWNkWKU1E1WNiope/p+IUuuAkBHTji
xeoZWBA1L8qM4unLCkz1kl7ewV1tc/KF/UA+NHzkCWFmV8wrSrGfWvTMuxKcpycrMUdTxRQKuTom
7LsK+nJVJ5VT4dgJrJScxk3wH+SRSg84j6aep6Y6knDzzr9eS+1seyyDCRD2dVUGqjB0SWge+ayk
z5fzsMISMfyufmf1MjVfFcZ7FXASuu7ffX0EvsO1J06QRggoDxMrHI69CFpHZA8aXmU1vB2naEDW
+G89GuS9VcPe+v+aiG+2VL155ocOUNCn7VCbzNd7N4SiztzceOP42h8cLtVX8+3BtRCvIUGj8GpF
L0tCuJXcXZDpcTRWI8uAav3rLdNmw7niA3S8fLL2bo9x+98YA4T1nQlw2qsDhkxuGM0y7GkjykVO
D8LNbhf/niLQtKZq4+DS22tuT++HmmnijvvFLGf1sV9uY/qe6H1ZoXAZq9C4MeCSKN/4Uru3uzb9
GvWRKxOqjBpx9K3+4b6Bcc3d1tusCHuqNYFFGF2G9+wMRC69c3TKi08e8JqZDQPXTM0CZhA2nr7Q
tK5Cet2gkyQUxDdPuPVGF8pL6ySluC7npOuRgWZ4QsH3pkf5RBURDouusBBuPEMNBGVjMdoieUZ4
NrNKi6Ztmy0ibl9TYor6ngGKCoH5P9IhihoUT9SEDUzlfWMuMUyU+0FOXOAwrt85nSFZVjw1QSnb
VF4OjV+H9ZMbxxKNhPcTdwJNqaSAu7jmBR+J04dGtbDLJT7ffsXoCh2Znereh/h2aVk+VH+pqM2X
5V2uXkMQK2m+XN+XbYVD+zwwzZ0EnxEQ6eJW+BFaGIhFWHrceN1rdp2HtCsdbDH1uToEAKF9GHvQ
ijjGTDVXIrDxdwRW2qq9VMHszmVDvdXsjS36SIL+J4HdK8MZKP5yeIMixlYawzstHBdpbB41qVWf
XwcxMBDH2Mi34ePmz9jWUZyJ1DFuhSTpeQb5d/owM6ffIrJoOiBVJesWI0gKBEIz2mKGWSn2smIp
/zzXVaxE7rCKHgV4KJH23o3GUz8aCg7BRYQnKba4gwy7OcMnZLUutDrn3dzdPCJiUZIRfZBfEumw
IYn+EAQHbYvWexgNmfQNmdcVlB+vjfvl+yyZIcrIhvHYmnjKSuzPpslACrH3ifF4BzMLVWM06/B7
gyroWUcdGhltwVauhDEEVhn19QyU7vslCGf0V2oo1KQgMTe9f+36D7QFZc3EcguMMg0Mm8gv8Rh7
4iJoE++6e3Sqg9kwrzkruculp719HXbH2E5MwHMxcoP1sLbbBCuwZpHRRHnpKmCLMKN/+2k19/5U
4tt2u6ZSaNA3BzSrZw1mPzP4+yzIBQx4R6dEh7JpMPf0im2TZNg1ZUBDXcdy3JtKsNQuj/QwnVrE
2s/pX9shqbagkAJ+TBphVZapKXcjutl37kL79h5+IzavdgQdB97HIgTy6yK12VMGiJg9+7HymM0r
QTsnTH7jP1LoS6ZZJ9GTBuTNOdvtcS4KftXGFgIDHMVwojzn0Guf+WW4YCYPFaszIx1wbnJ5ccJl
oWH9Cx9zVgd8BTlsW/Oc2APqM6sTAwc4RDd5j1PVy4d7DIWjNIJcwLx3XedCXHyTjC5YNf4L3Fyk
m5vKLxclJ8JwDssb9Lw472Y33RDo7gJ0TeiLrC1vajLYuspYGlaHAxX+jZh6Jf8VRBsJ50YXiBAo
eQXuT9Acklpix8J9NuVcTmCmjK/eTBa7diAVwEhA5oPw2lZ9yB50w5oQ8MDa0MwShGLzL05h4QBP
GO1GGwBFmV6ikazxZ2GvwK3CbFHNq9l2RRHpgvU1/cgvSEIL4nW/Nr6OlJ5o1XMoqjMvRz078CR7
LCIWmIU9coB6N4wHBI3qpuiRtaqK3Q6Td2CgTHW69IuGj0eVe8sjkqci+Tc+cyas7aY/WxiG55WP
rQPrupd954QmOHJ+4/N3FmKNLa7KiyYWadnXXFlNG4g6hiZBPbVT46KwPo5nmC+mUmwArwC9Uoug
hAtbD1345m+LuIFk1uz0dMZnXGd17FdzWQmuAleX+m1TK6wkRoaR8we7Rb6pAp+YMQjHr7ueO6Mp
wOQQD8HglFg/Gpjr8NAlC1jR+hCJw5pOTnIt8xMJyqOGv4/AOq1iMIB+f1fHS4i1+6ngYiIDRcty
tw+Fhe9sAaXECoV1AWWU+92DEKJ+sAkffG2//H4+utev/UVjZlH0N/aPBpHATxW1cnUrctOsWjVR
yheD33aeXBTbpYfHzs3WlrHxXNeEEMKSG0RiSOYX2n9GirIlmFNMDPpS+rYLghSXED9ibc8d0vDM
WbTPpRn8HKVYjYvw/7n+kGUQupyMU9OaU7sb9hbWqRKF5gXgaCawyz4GcjrfXsqTTnZB/4fP31i0
+OpZDKOObwtJHugkeAHXlsn/9Ry7Yu7xHRfhevKeSym90gx3mz5GdC3CMMfpOZqT1OZkCOt7cQcf
gwCbXBWtie2oWr3dMdp9j7Yyag+PT9E2GQlsLk0xbF3pjSoDP3i+b8m9WlQ9oIuuxRc85tcCilS9
3PImUXtawEKwgk3s+EpaxKfd+9l+/hovTJm/3CfU8qH3DBbcphwxeAlzqj5Md9hxlAMzLPpVPPwn
qcRbNIgeoYMrly1Pre9dNjRfwvlKbA8j8iIV1ENR34MKD6EGPHrIc9MnokGOD0AwajX1ra8Lrdml
6r+nKTfAPtgSBvDO9y4dgwv4ZeSOklZewTy4tBh1/yUsJ4XbX/qEIkLWzsNU7E5jFQud0tuUvYTc
cRlmPdgf1VoJuQ3OwYBAKjEovVce06HdYRTDC/SHkDMnHvQiqs7fTQqvr+piv7WVUvrtlfI4IjHW
xtJM0p3fDs/G4hhvP25qhbieg9BB1LsRTk4i3WqYllmYAkS2MI1cgKsD+n++6NK/mIK6CUstrTrn
m+WJLFCmA80r9p6sCsKWdzkn1OOPjZXg5dda8sydzXpl1CdmlV1GfWLsEUp0Jr6ezM3U79s6oQpu
5LJ7gdmCTu/y8L4pZjeIJ0RxARDcEYHzDg0chuGrJB6TeAWDSjMe3fAaqtlwj2bC0E+3F6/aVQy7
qbW9yU8sCcv+mG3SQXnCCgDkVef9v+0M87lG139L9PmbE4R8rieqDIWZL+fL8qc5Sc96BBQYzIyM
MVGSzYtYZPlw8tDtHaXUY4w5f+VqvRTSjO2RORzve4aUxfeHnwNKglpZrvmzrWOJmOkDrRA52+FB
jCH97AM4/1xuPTXCjlc91ka5bTDlQlX9QUJoWJ5LOSRX76FHebtuCcDlug00bBn8hfjg3A4hauOb
Orm8RwdpvHZGESkkRZrOPLD25UXqGNMGdp8PwjwgGPi5pONdAuo93TWwisyfgwLttXOKcK8Vwg2h
p7LwMcLNT2H4ZeM/i1ovwx2ZrgCfb1brz2r6E+JLe+luL84mnNnROcBpsLygmhOHfv0H1+PzI2hI
FeeLo2PYNawUpxgqcGoKhEodCykRWqLmZKnhazbO4fvV8UWTBUevBR/Hn62hjJtedh2IH9r46k+u
JnBh84RxLYKhRkc1+1wL/fypdPrEDqictOq7NPtkzCAi3ftFYS4mq3eaZqAZAm5ZKxpZAqvUmg2Y
enHdxkUinLohMQSXSTQd2qfW1QoC8Kx/XfPgwx2dIieSf5HmFcHw+SHcKW8F1IYMbIkvMv2hD/h/
zgRLOh32TorC4rvjZ/6YIdEz8auy7ipc5/qUoToongujcQwlWoTm732bFupGzUOB1kHSBF9B2e+E
ANz8uLBxMN2csttMsKHLkCw9/WM0vg+fJZCcJZkwlG7WZ1JL3MKeypjir+igBqeRlbShx9Tv8OJm
lo56mWonXPnHZlT2K55nd9pw7S506GFxxSlrhkFOXnv6WKpxUhHjpcjUiiXVnGsznwLls/5/4YUl
GxOfNK8QCmvSTsgGLEiEXP85IZSnJ+cjeXdvrIvp6sn+n0otJQGsRt843J0vUHkeDcM7X+7KM/P3
V4HyJIWamnL6lq9ZnN/Gb7ULkseIFhU3icXZIwqfYZWQb8okTmQNhvzb6kpoJHxonL1XO0a2mqjQ
WwfSCd+LynfEu1jPPLWUBImXLsI0cLhSOGcm65YOiNfbAkPKxOknRecfzIEI28ktzshN+WJ0eMFf
DMyj8iwNOiiNKAHAwr42udOIJ+jOmYp+so+Pg1pyh7JNre24yokNE8K93sdgOrs2nbxXmHoZQqjm
8RxonPJwTI7dBOrBjh40HoSbL3iJ8x/HP8btxtCPWoeMcKCIKsl1ekc39AEAgFrC1/PqVbit/uw0
kRWH6ju1QznfyzrycaxcN6j/F60VWjA8rBIZ2iCwGm0c68wOHb05vVzxhCraATR3D59uSM+Nm4nT
3vQiISwJt7HtSM9yR3UpjdWWDp4eJOH4vBAtBurFkdr36joOZpj23RGGfdP1Y/hiF22/foWp8rdc
7Bp/ZmMacA3udJb79BTsC8cJ282M57DHcsXvbTa6FeV7102AH8m+eaD/YKqTXTGKVzgRchosUUfw
RrtXaYaF/rjzxLIwhxXrVIvUYs1wiskdhB2PLM6UpkR8W2Ve6BB8dZEyoy3uW+wM6KvJb3CagNM/
SGdupq9siPJqcq9ZLo1kLNWTNn0MQ04q5zaZo021qz4m1+zrNb4SDjc5VYe7YTDEKePKOB6fbiib
M4W1C0kitYk7YPMSxss2wnzKt4n3eaeY6SuZPf4YELvcLwpWdG57hFPSTcg3y92Dkv909DENm8yp
s1NyAUvENSO8mqnycv1wSW38DMNJaL87gNDUkP4G/Soyp8eqPdLPgh3IIjP/aek6FbtHMEM3vHBl
w0maZaQQQPQ4bILXM/tPkLXocl/RvANoPZH96zA+bCVC+BBtYblA+zgL7K/F+dbvGjnpzoViRjoB
5XE2TW/ILb4QgN8+rIyOm0Dhtx1n76jCP2Dk6Elu9LbCeT7BzL4BwCi19cFNamtjZ+SvpTIrOy9N
acD4NEsnFqKeP0+jQgVZL04+VdZQanWYiOgOljppgX4mh020lF4b5a05CPbmhjffBYoPztYagntp
eyS6UbKG/N1WxzBSgVVJj5aV7O01sFJMHmw+rXpHvvyF7pqF4TIeJSv38PtjStIeGa6149uyBAtw
i1sW+o7fyszZSDInx7+GhQAbleJnYXJGaH+HD7+ZSICCC24eGBj9TyiPGyf8TtjjwElDjFBGhYzK
KDi49XPQbd11B/sLdyCVOVy3b2IembTgw+R5mPYnCI2HpIRO/ffF5tfw1tppHgQkiZZ86dzDsA3K
Q5pUAK5eDew9lHwjxyC4keAiAf9IW5sbUP6Qq42vOgCDmBFaGSNlF7UnONcgJHYn/W5Rb9ZnEPKM
b+WZPnNW+ZBp0jtx/PFbiyyTvCTioCAAJsPrL4BwcO3/bGHMTYx1t/aPQAs6zreCnRgh3j8wMMZQ
ethIafo7BWXwD4xXjVBvSNKAFiJILTmBXhcyF1H8gt2O3eW1inadp8EFqOAU5Z+BHQUovqeq2JUC
GhT0Z1hEemEmdp8BvkXLHP9MVI1joSJGuUMLcuV8pcX6rg/I9xxSs8zNtxHEc/QgHaergICGvrH7
Zlc6JSywIVYRM5ETqkuRzaIfW7NQka30UJXmksEaEtk+g0zpDUnYglJmMZgXcTOM/v5NEiwgRoHg
/watQnz6HIM6/JC9mVxVbIOYg5rZ2HB4vWaHwGfP5hc/g1BBqBdoMsmvaneL+v5LfCTf/WW+/5H6
IFKM+bc3VJ0HPhohgrY3VMLGDEDBM1Ry1M2768LUR19aQGs8YYCtOeMGZzSi11wGZJsNG3XKj74u
CacjjAF1TL5LeTjj+QJDVBG0udwsyX+OfZTgfIPDvV3Mokpl3UIPCxbFTbnOqwDf9CSQqeo1K9hs
C7W2rrf0XV7Mgrc5ZRdRbb+RBqaCPGUoOKR0/ykEwxouNhzxvkFgwg/WtTrljmVewPYm2CubrVku
KUaDQEtfGpXBgDFJNpvzwS+fXLqb2c0bHtkVpURDlX6wj6nPd8ThOZlaBlMgWiRk+j3sbqOCykGX
BmYa6skBK3L7xiFLB91TgjPUGOWCz4vvt9VPnbWYANWMRFriAecAGgx1z0rHzEjMBHs/GYtpfzti
DeIveUn2aKOos6ZtxGDdzlcZXLZzntbVVnOFtN3NuDcjyeAmJHRywsuqEfqw7jVEVl3h/ZUv5+3y
Y++9xa3BSNDOM3TXBkZb+uNyNQ3YRMTbcukcHwzl+tt9g0XigDSHabkaUbhDdFii2d4dFXEotXBm
+QW7AJwBgTK5XUgz6/lbozAXOyuuuNvy687599eXNbDPB0nGy2+EPmYjjH+Q8TNQhxwFBz9HiPuu
7zw3lZlfebS82oYQKaNb54lDyQ5tlaekNOJ8K/VuCZtVIcsNzdbSnPiXSjkgtP5rk8VpMjRd8SJU
25nwdaC1dGmoOs/6+CcmMrOzxx1xedxWgV7qxuSmj7upSOD6DwvShNOhnubkGqGlxeQYNcYkTwR7
IR0lbHbcIm8qEKCH3ssJctgztqokfBmnVWmjVb7kWjDcyaYtEgkYqyBZc2zXY8ZPPP0FT0e3uMqp
sFbmWT8+fwKkWoejuwjOiPGJhiWWh5g0YUU8WuNENN5ZDi353i8az5JMTeihuMDALIGFRLQH7Fkd
CBhbeYwgKL2BLNOh9EdfIPI1eXJ861jUy88KM0wz/RyjiR6JWB7XS7Iq9UmJTrHpNXUpahihBpja
xGTo6bvjjVk2EiPRpXXxIiMlvJuNTqKLXp8KNA4ikWBxd4BkDkuqLWRxKBSEy6XY1yHZ9NKkqY3w
gccMofKa3afEZ6J3cjI4t34ivAtQpqX/jjT+RU84jR678mEmij9TIVSx3+4rp2kkwRTueiyXmIk3
uUvgtBwvIBC8uRRahuJzZ2BgGv/4gwU7HM/oW2MGFneVIAD2i6Zat02mxNkZ7k1EZpfHd1cKlMg8
SaF+XxEx5uYvpwWGWx8gFf24Nv4RcdD4AqDYQ5fBdNhQAVW49S6g8u++LXullNSdBstb5OYAZikt
2bgsC8zKBDpepWdRJu2DSZccfaJsEj/9gcnOUghfwd8LNtN1DqEkXumJR/5x7fEKMw6FPbKr9KPd
SakunlleWePz4u28xg8qzrdUCM+UZ1s4RrEaiUi8xNDHfGOpQyEsbPqqhnvbE3On8UoW88oKhMaI
RqOAkPB+PCKe3L79/Juntv9kx527UzgJHSTKzRJpEwrIDAPwTht5F8+yiNGBYkXuNdQJOLqFvbpF
GfH7g9c+IJds42uMnGXcUNPua0IR2fqtklg9uvheWcDC+1Yt89vyhgaVWgMTmybhmI4mhJVsOSts
QSLRN0sIFZVMTpDXKZ/hhUZRP/NSH7ITJZFy/4rdPGLkmFsFOTVegbIBTkXmo8sunEn8fsABdXye
kWqhe8+gxnLr7b/lWFK5z/nWEQC+FD6GGJypYJT2xJ/+17BktsdT+bNZHYzMLk+JS4zAKoXX3J6B
X6vAAPYGvLld03R5y+8pAN6ZAafF7OzbQgGHDMkFKLFV7t7SBsnMXEO5QdbTtXTpmArtReDeCyRo
hR6QEABYuUwQhASmy64toS6UTA01urMJTwJzXf+0zy1zm8WMg7o0PaxdVnNe7MzAOhfXEIMSvcRV
ooW+3qbWTraGOGcEwR+/jLHwkuK/vOPPryRLKTDx9fmH8mqXsA82LtdCESxvTuq6qZK9NVn5iuXs
i3zOMkffmECWLVSaR5F2Er8A3Uy0QGg+ixS6UBtPkLxXS5SkIXOdm1c0NI0QQk6J97zNUybOslv7
Q42gHgiBLzVMJ318Im0q2VZqeJry2NjWvK/JStoJseaPONtp7Z1t3did1BvitbH5ipOgkhzoBtie
ewLnM21Ja5uUT3xQd1kShH1UynesmnexT4jicXHMkr/HmyCvMHt5ax4AkBhQaOu9Rrblk3Klwv5g
jh4GcpDuyku85BDOVvr4lTXqkXZLYg7pR4XAcckoru/fTVFmIF6cKF3H6KceQ4yoMueEFQLOyGwW
6BKBvz7HfG48QpFa30besvTva23H6FsbcVi+2Gi+viB2YLYidppMr1DabE+v8nd3478eEuXZa6bi
BcOTw6wBKDh8asrt1R8mph5y8wJmWnAAvXZx6orpwJvY30GqH+ysrTL+Lh/LNCQ9+Q5UnMqVFWVV
lqsnLOIg9H6gtVJ18ICF2A3E1otjV1BcdgUt/WLviwlIevBM9Py7W9hnEn66lC8ZG8zfXCkPWw4N
fRZv4Xwf9onqSaqKQtlnIjLQWLVLRYEh94A2Mjo/Xc5iuMjsYYtpAlNdpwg/aPBB62flUM3JeWPh
hLnywxLuIDR7TyupU3Y5ZbHu1Mnkh4k1MyKz45b+zOwwBu4FmFjGXLLSn8f2EYMrqKqGFs9ytguR
dwlIC+wCuKXEbjPXrZoGFPjLpOprr6LaDvjsxJQGBBqk+3vQUBGgx0KqiG+y1q+GEQSWNrfJlH22
8c3HPvRayYHmpOngnnHM0ewvHxRG/BUmzFGse/CQ6tHUPkOa35Npm8NT+AZWgUu/Y5f0Ky9pGivL
Q/JrGEk2CqiWvW58/cjG7GuG6DRfG4FLGbx5DcEtXiyfULZcdFUxv8yE3cKGUJ2BKXPwaY/Led3R
mf/8kGNjex3xxkUAtIpDNiJngpSgHkhlMESd/mUdW6fspdTfCwY1CXycCeF4EDzBMmy1Sim+POuB
jMXRpmhOPhgofdDMS5kCJiKxawd43nr+lZamP64I3GcEKaXa4vqzPmlYT0NnmoxWSpYMyM5Fu7zE
dpamnDMAxscv1dKJHCI5UCb+7Z6s4aIdgG9p8h5ttIg4s8qY5HYXQ2ab0G/378ubXt4r7W3FM+Qa
daBFDwmSPd2TJwBXFeE7jLb12P6yIcYhIwbbLKgzlBsrVdCm0z+ZvLUEU2U9D9F7uWvo7xRCnBDY
Qo1vx4f2/Ks6Gbm4ZdzM40CP6cLsFK1k5Gec5dyU9ozOhw9Z4znFsCfHYIC+YNGWwPoQwSp5uIw9
ZxhcowjahabnPDzliCH1q4o72jDXur8j5zhUZICY+uaVLl5BFsh1PCO2BD5BmWF0psPZc+SJ5cgY
nWgtaAXOHn4Dv76zgVK2RCLdmB9ZDsTffvEuIjXG+/hpvApRjBMU4IbDRFoA47KOxNLttiefk7+l
nex/7hPRewQCT23SUACsTyD3vIRedqMpG9TO14ZYZ82Riog9fsWAOo8J2mPUTPaWKgO9BmgQeYdl
CrokZeOmIXc9/rB7DYXLR+nRqjLmgCcS0FyYIaLrIyNftcY3FO8Ef2bQg8JuPm+DUdrncucoPHOr
+35N+ifugvSG6iezJKPfV65yvCtSf3Dfg6qpy9GhaCCHJLMRqBfn6+GSgQW8W3JDEH81igdEwjA8
UDfNTU+hBtKiQwUnbLTrszOS1oFlVZM1+XjgmCLYfXLQYTOFE0+V4NPYSfhJJts4WuFqBkrVQpOt
QXKgMvFbHlUH66gVHelFrwtdw07n9sKgoUg3xWxMYx1Tc52lXriLnBmuacLWJH1Q13erv0YtQJBO
zs7vwePcTU1P1I+tNeTDPjKxjspJFxqjxma1moR2q7Jh06Dg+q37XdcqyuktO4gXwBfnTELSeiYr
Jv5LrhlZyb6gyDY1a4MeKVHqlK8jDRZHUlvU2JFZX2ahcci7deDq+4aMpwjnrhMgVsXoaqZHg0Zt
HIJILwNFp/jfdurlrKMg2dsL4oxRIGU/5AckoDpBOKrOV+OhIT3nfO4r4PwLU4FXuwWOEtc772VQ
rZGdyT0FZNICZiSaWBfcpvKUiCfIVoT40f3QSRLvYIn85mjlKq/7k3YqUbLtNDcUcUfVr9rdylfK
6nBvEkm6Cgbh3sQlRgzZiVW3xVr5N2fvAknHjveyr/2UqHNMbnHDi5kOSe8seYH5T69s91H3Mcsw
aISfoFKfiAS/xlW8/mykPn1TqIaz31bDlL6D1aLQnj7w0RPbkD7qJ1563CpbNniSBx2apD9jrz5h
UyQXwqRiGGfqLdOifFNjfJCIn8stgKs83AFFuPxfrNK+SurF5Cvixy6Hl13tt+7ASFdy38xqjCav
mipESwOfzDWbM3IIiNqOsqeUFlG0y0493oeAhDMe2ctGJQIrswdCpu/YQqmteI+VvbaotiJ5qWNn
Ey52Ql+vCGl1By+uSGHBMFuUA8BVYA60rT3gnr7MVxkgiMVDrJa52JoHcQIaRj2CEHmyTm3kkg3l
JQw8bZhRfseUnoj6NkcuLbKRhcA7IOb320dq644J70FmeoAkE/cNcLZ1oSNQfHSRLQ9LJ3Wip5IK
Qgvlu96nck1FdooEdb+yTHK7HDa8/L+19CG96NXH9LhE5ivi6CwTg+qr7D0e9WYY7y5VE0n4SvOH
l6XkMbF+CVrBUugh2Xtdjq/Y4EbczBFObvuw/DTL5lYrK6dbouZabl8lhM55JZsOqoMybJR7jB2s
Bte05l1GJlsupWcMhJ/iXKDZ27s2sh9QQlkTCPrFoLNkmQV18EznephabN9x9rrdJ1agrnj4bZCn
IpRy8SNCJN14x9DzpQHHY1zliuioDT5Ow3GZhDhqkKd9s1QAXQtYHiiLccmDL1XcwWPW/M+RxwsD
+uRnQPljcNrkB+GCS2owGhDg5kCpIpLA99VQJsUihY5XAynC0E8sstdlkWmECH/VlTdjhoTz7B2v
CHmqJBMsm10PwcyR4sZwhT0W2ynKxOzWbpGY+EN3LT3a+oM94acNZspguY5UYappoEMmOPtsyygQ
Oqv5XFRnaedb9qRcUmp6O7ej026N77SbXlqXIM1kG39b2akHojdUf9d1VET8MfVhXLXINd5W/chK
LdNEdX6y+Z+U+I+BLLHEmsMC1yEWH/zpkYOfnmUaozazQcC//jcBiQGGPW745sY4sZ4trnNfEmt8
3H2B/yZdyEF/Z6I5Cda7+p5BgB8F0aPc7KZp6L2KtVsiLlKPzRnUAtR2lB8QhhPH4Zdf6IXA+MWv
hSvByfXgzHofgJFVgH7shoX9F+Pzx0qDYoVoeMyRJGeubZpAv1mwCUWp4EqwNtq61z9Y6u/7eMAD
+dRYj3EYQpn2emqKbBAnc8eq++b4dFobwYQ9TRKDUiHu/1gyntT5Mp39NIl5FNOQRy6PxF7KcnmZ
uOk+ltlpq8P6McmO4yArsJFpRQjnSfLVJQEBn33UbPs4DeL7loRugLdJMNLBaXRIhqxEyv3NMQ+l
Qo1upXhS7cNccA64mO+1zc09dcCqc4I7pMzsiJCrg8Xm80DQ3o7JP+ero+bAb9sJabDo/Z2fvE43
Uc9+u3Klpl6CuGelsPRCFeVLF1vFEcUxs+I9n/cxbbV1X8fZigAH+H5GrRn5w8w00WG+bZis240q
ly6sLmx4p5epBPD0aMO5C8XAINm/1kuSq2ZgD8tYYXreM1bna9BP9OLvHY2Tg76z9n1EID0j5jOO
C2Ev8svJxhV1KQahkFme7gmbsvVbKBk6kK88NafOTx0nd/6v1NhPUCQSuFafhDcuDJm4QsDyix8l
HYnve610IyCTyPOgYtr1gFO4GOsIsvcYmdZHgjHeS6oACGf/8K8pBSGsCcnh+3Ib/e8O+hRL/zkS
hr1ohfM2o+y3EVDn5TNqrJ6DpzO9/Q26S6ApqID6VDO06mHA2GHlJMLdqBIWoE3fcP2xPXmDkXi8
HuJ69070aTqloU1HwmWa//GeeexVQmmgafMMo9f6OEc8vHIgYk5en3ONGN/dW6RnNbuD4yKnr7RJ
to3yltr4W+xfF0sLLsKb72jfk6GsRBwsENjvQUaUxtrkVreV0P5P8A9kWY50Nc+S/mtpUUvjM4bR
tjO0lCd+un8urG0mP+RaqjLhsr/joX6ge3OrlRslTmDov5kewK1Lkbj2QO4tJrERWUAgfO1qIfsE
vFplezSG5V4RfQ12W5yE/A1Tp9BTM04OkGk66kC5BPwQiIrO9YtHIjqSBlqNiMpaTniD6z1xyI0m
6+BjwxqrH004N+fKy+g0MMSyMDhqx9r5O7Gj7J4QeSPza4JFbNosoZf47QtpJcOnjXI4e71Z9gMI
ieXU0iaPj3u5LAa5EV8k14eszhOLhP8xEszVQojmjbku+mcfGD+MtRJCVZbWEIqCmlBYpoRvmXTo
xa5RBi6fLvUUWjDrGHxNpVjlSe+6dFadtvRVxEb+AbpZtyyUScLwggOiZ3W/4Jk3DJcacvSZlGg/
B9iD/wFZkNP5ySBpKuj6wsrVtATmPJy1GqUoaMW+J4iKOzqJoUIaGvhXUmxK4FEcX7jWszvyXNWN
u+iuVR4za8yAKRj8fAwwNZAmS8Y97WHQjZ82CexzHE8ubd624DwyH0oQYTY2/XfiWYU89ablxmIu
zyxCVcyfbK35x5JBJ0aoe6PXGBRHY7c+UHgl6DjJ9LQDNUI8Dk2ISY0JCR+WS21Bf9s5jL8S1j3B
2diFfCbDlzMJYUm3BmReAzHc7kd4inRZCGsJlmkVYogLzjXasKnFazLotjPfrm7Hasks/mSMjEbP
MHDJCoR9fIcBjDCCYlSLCYKASgH+HBiIbr+2iNWpYAaGyOlZupTpvm65bDoXTsZgW9SvcaA+gT7z
V2w+RyNw8Hpcxlz/0n1/LH7nMOs5WLNlkrZCGnAOCp9KDDYJjkbSO6eZyIqvKSFZI9AE/8yTRP6w
PNVR+jijORTtWiL999nvdyKiDyJ00n1HxgeHOoBYQXMNvzL2fCK6QZ5mMfmt26rg/8jPWjQgshSU
vRJO5Hl771Fbf+nyNoGDG5SXgvM8mlQQApAHzWnZQ8FIWc9XrxBnVh71l88UKX7gcXCSKBvHym1i
OEPBDdocNCedNvTdnZoD7ANmEGsOAXuFc7/x6YYuwCgoptK6u3zSeXH9HL4aAOautQceL5EvNNie
8cvXfGHDT64oaHJNUbMXqoDUJjX2azxuKkS//URNvOa22IiX+KAya4n44aUjlxv7rpy4IT1ihwnT
a6wygAxG3ADMOfnL9PWELZCSJqLPQA/n/MleMJnHlOzZKLU+l/CjQOTw2ya+rRLDKpq5Zko8cw8z
36MCseva5WB/h93zIu1FayX+3hsOG7wZhON6LFRYRGdkVOwmJO6e6QMVNwvRlVjA2VItUri3rqzG
4GgsKIXhwtLkyFDSZtmBq0hweJduaMpYoO1syIeXkrCaX26vbYzvIe9o4ENa+QLM8Z3I8sr9d88G
hsT6bWnLxdnjgfq/Pj3IvMK3MvNoyvzkSkFlP+l/ziLiQRIO+26koSBq3wgxXAwgynVJypkHBXTu
Vw6I1L1poREXSeO1bBdLHQC6Xf3cDE3ZSfIZVeAUA1vC4DBYNxjYvbqER4dD1AfO1VnJP3Pra+eh
3/raq4CFfD2dZjAjkRpALROncY+7MwQ7OoXakwaczV3yj+jx/ZiwoxQaNPJMN1BzOHfUxsEM1uFP
TVYsrzDn6KxK26Caes9aUOLv4Zd41l/hcbHHqq+rgZ7MjJbBPGxwF49X+TgKfhIzywi+69kKXPMi
1gam7ik61ceyf8WLBj2YH9KGN1cEThUIkWUjrGp8217rtgst7G8d3U5KJlSQHmJnHmEaSboqM2eh
b5iUHTBQzbrEIYQ51vfVWOTVmCgit5r6HkRufIIuJnu2MKeGCutGJbzKQrz/JVT53IEB1sG3ceTJ
R3lZshONIMs5dJMRolB3d/TZwyf+4IPQB+kQNjigCFi2BVC8IqQ36LlQ6LpWI7m5EGOWMLHwdQwF
37lxYi/pTSiMY6eoEBz5CuO/TdNvspIAMk3AQGTlzwxQvlVQn9P/l/heuufFi9Lt+xtUfxvkruXB
+SN7tJc13S52KsUnTDNnZp82YYv6VWFODMpW+v+boaagBvK3SXj1U5D+pw9Ozy3Q28qthVxA93/G
P9GzgNTeU6sCiy60+9O+Qua6YqIvGHWxOwfmuN6GSJinykj/ZSvY7uWTo8QBkcJzWgUEhQMofWbG
DgqIuW6wdBmOhCGiSsbZtsLfFWqkmEK4YIhp98jwlP0jCilpczuJCdJ4EKArf7P3rp0oR4j+/BBW
pZp/TgEXBTXPVEeX+anbNqY3qG14QwoH2EbYwCGF4dFpEr1hrjm3Al4+LGKiCGc0gEPRuV4T/Wfg
LfajA7SB8+nJXPsqrfkFZBZTyUmLQIeFN4jk8XWLqQbvr/9oSki86xbJFGYt7yJOwLK1jUK73mJ4
98zjrbtWFrDxxu3JAk/VsyBzTAtVefmS4B3LMQWJOo8BAL78hwrh4SnoSaFioxfd5b1dNdeB1bK6
B3mZ9H8/BSxoq/TFntivB0qxQY8JVLATWCryPLesLWDArB2clDxGzgktNKAD04+En/F2G5tHsQeJ
l2o9Hbb/EvdFVaQWhT4axnYoFejEuwQrmNABO1GZPMD9e+iGxLLSeQuk+Vq03KLLBwUBLcyNR9Dq
Wc9VgFtzYpcZhilxD0m9cVdavZMAF4MJJT37tAWXsuPyViLsXdJEYvrEqqc17XJp1OvmbPlyRL4b
EzQZ3hywo1BLvusA4VQ+EczBPrQU0PwQG9gBTBFcovr5QemPcB4l0gi3bERkdIzbv4MRYQizSkSw
QSq109/MV1VnuS4YvqrZL3Mi3oTql08eS5+TfeAaOxSXgy6173WzJoMhfFBplC6KWzWPY3df7J+k
gKlZWgnmCbcELPXhM6ARhvhbk6IuJVzHgkr9KO4OgE4PqWK1ogeg4fWz8H3ZNFfuC07/f71KVfjY
wcR/mwKEca3H0dVziOYZnnR/BWK8o66lsaq/f8n8hmFctlagDKJtbqzOBo18UaVyowsIygBl3XBh
5nBErUQX0VwarEyF88Qf8MTMBqfmWprqUD6oP7efRnci66mh7gayMG/ln9pb/SfJKR0ToRyf2S34
wL4J7npayeO8OWctoVtCRPkyI8GAEEVygBHmIqIQ/jgQjvM2sBSbwy3lIYgGBXhF5ucK6h61B5tU
0u2esbxPFanjfO9oixER34L7RkneZ4GO3CEBjt/N383+TC95Z38lvNEvL56/uXka/gNctk+j0vzu
PeZOkmEK9Yvoem6mSnk5erVeieY7TWn+5KWc44sdzaJOrsxV9PidggJ/8JX08GfjFKrgq9N5qPnr
E3VNKFqjZ0PEIDxAK+Z2OlGTssPbTx+N/MQC2bNzlURa7xzKYraurWWJL+VvVJnGn+E8PU4FodbF
LEM5bOSeud1sG/fLNHvHKB2dwTK/LrRiHv72EpOX8D2GYdLqqtsKel9RWW5NIX0f4jsMra8GYya9
2EKCcgdiHhIVyF0itgpAkwDkzdqcLBNgY570/mq5JKR3A5yzABXqAiscAh5jLl24pWB//cqv5Vkm
0AyEIIu+6/s2W3U8XD6CRPbRBxB48Nb1ntR/xOuYEOy8TkN3PF9b1+h+iDyYkjnQGaF9tJmkE8As
gIt7f8ALeWaNJLlWuL9pfJUYX3BrfLg5CtzCWhgq7jksTqzTcs0NepIr8TO4r4PZpHixiyf9EYzd
z4LaAyuEZrtyQM7PQNrGB9h0gQR1dQ6WbPy2WRdqy5hRb5tJi0TkajgmGgt2ddlXsPEIsd9oKAHI
0YDBkg4wJwoOIWh8fzuC7mN4SiaKccUlo0oLx1AMz3uy9+yEVFmnNgNPFiriSXx/avlKM4HTFhWj
uNPP8zK2e2fxyHbGkolVs+1LdtveaaXyTBveTMRvohu5hs2AxD8ZWgkK3vRFg6G/BiEd5MBkol7R
UrkovhoodDhQsFi26J9yXSoNoPKyFWJ7agawc7isdGh7LRrqxu7uLucy5ermd33M8TdJ/+vIG238
AAV/buFdr7g3Tq4//2WyFe7ezpem09xr45re9a0HYkC5/4HeZxD2ehYG8yEZgzBL+Ko7aPQmCIik
tje/7iyJCjCZz1get/JA6JY8ahmCLdxo2Dxi2dJYctQcoMLBgwNNiFMqDQiHNDxXLe+PBewRlkPt
Ok0CeMxSUdOy98H5Hg5aO0hM5QG5OG1u8bs1xHWNzDUTKIEurKKgu/q9zzXhk4XqSMqxcTdcIlUb
1RfdQladSvugukufjajdgf896bjMmah1X321AWtlrUWlPCGrGntEaK5ld7MOyhOEGDMiGydg+45y
VOCk5x7laseXV3gf0EKBJPNLBQ+zA71fMa1ASq2AaAzrCP100pufwcceq04HOFUe0pyqya8864ij
QuFiOXibP3x+2hGCurdRZQ6rty1IB85F2Ykxu112Y87szFr022bH4q62XZkYW2FqDXyyI3Zd03cX
SFJ+T8M7A3xvdXcPW3Nshvf1/bv+2SYbcha8r9i2GwTfq2M/1EyHO9uMyaeCxFMYZYNAOL61PAKm
mrk6Q13+lhIWecXgMb77MlHIh/DJNwTVHcEhQEQIhLXLC0L99uxvX5sSGJ6MTY2y+2ZiIMpw24M9
kumZU1FAlRCmGgjKcFd8eN0wKS72MjGyIflKyqI7DzXpWvjpEIQtGDCBhlBijyObZI0vauPQUNle
+UwfeFcnU9ADtR8MgcikJyBJSA24ifAHkFNWhpjl8yEUGKrtXgCk0U0cyVmcbH3ThI6QXtWtDYzO
QI1F1xWR+15yLK5ivb/1bsy5vEpqzIc/R9qysshKYzpc5nwD2sxDOvMVkhMfzQ7gNQEgSshc3QqZ
Qj3LOTklvKxD/D4sFy1ko9UjK8YxTuPKrVK7bm6VPPW3huf4+vaJv6/SwDrp7B8TURRoKXUhHsJ3
Bae1cCqZ5UNRtj9ps8EEMSNFoZ+w3UnyVpTGVIytuW2CaEZ8EvnBNfmfsRHqFkTxFVkVWhtHPb6b
n7AY5aBrPCoRmq7Sj2KCZyeCnCsiC9tbB/hiSvG0TXVACcUW8qg8lnAb17rqA/sV0tQAJeEBE+Xw
ZS3hk2Wa2TuytOiCnRTFirMt0KAo3ygvkC4OzrWb9kMxb/H793CnEMT81JQL9hVbFREbAdXVfFBl
cs8HtVG4BaGrENPo215Vk9k9qGoEefgyt6MTzmJpP94WoMuffEDicK6YrjmTWBGWMSZPZt4gk+am
vDiGGwfyOkKrpkq6Xop2L5SLgBcXpPzmJDPuz168ADltF/krCbZqB8Dup+CpUt6XTAez0m6ZIvDu
xWkWAWLjcopVAtsrtgao6/HTPaiiYzt89h/y54xdNCQmyGKdPIicB9GmAIgOhCrSAve7QGJuYG8w
25IQxPO97Skw4uH/grs6I8rFHz/ZRtsnTWoQ7B7JEDwBWbrCVqGIw3R6k2ltxDm0rWynMH5kF/C8
khbC1KtHd5Q2WVlZUS997uWmmELQH1TALSO9fDc0QD6kT3vBdW1HBtxrwR09Abo4I8nY2qU2B2/F
dz8/VbsYSUlRLZknTJV3osJBubiqWJO1y0DZ6Zb05UOmEO4h8XqILv8rUb3k9FmF/ebAI2A5/YOr
Se9BNtLg6f9kf1cKNOo++25l9L3K7yhagZXJQXCCR2UblLbnWF/pgv56HcMd9MA2yQVnt2Poup1Q
XBLQ4FDa15j5gc83TWHUftfcUlHr7iQhATcBCv2KHpUjdQX/oIXcOqbw0GenJoVl6gJAJ144EGuA
rM96pNzt8bg1+aeVe5MGbG4IxIkEJFcraPWQ2F1M8SAKRSYjg4EI0sckoFDXJd3WE7bWv2lEF4oZ
6HAdvxDOxVR4TSmpdFf9IrtbDy8qYL6pblmNZykUmdhyUkz26rx4LsjCJx3mksCh62weyo9OKsfs
M3zWdgSJCEdzqTyDjIFvk46f676Bz2x7+YL2OXUPVqnFAm+CrkoLN2ds5rldgLTaRugNkeHmTmOG
ZZqqozbGpxTrvtE/YN5Q39Ike71xm4WhDt+QyRU8CFTgfOEaU+nTGaQOMGHVorYCC/gYmHZ7ZXpz
JHXYWYh8e/fkyfMj64IKg7oBtTU1ujn94MYTkzVVh070zSKAMlQI2HJxMxLtW+WUZgNJlaP7NTUI
BWWjVMYY8yc0kRsxXtM3MfewZzDAzRmnqCSB5HGLu/3H71SKYBeEvQvRXHVyHxeUUFR2vycTxL0g
qWeT4cFElpUjRJH+iS6xvxcwOjA2uMkcp0kKM1wK1p8Eo3mkWU1Ha+mj5uor6MSIjZ8TJ7tDQbT0
9779bN3XVciILeprQJYNlWazDUeog5S2q3u4hTPuE3kKSoPIDGeYUe/gsgtN8+R/FdimbJ9+93Q0
ZYC33RSSk9VamTpwe1KPShW75VAtMU8iVml1XeE7mMYHDoMDLLVoayolZR02gHK64rXNf6eBcOMG
ivhr3coetJKXNvIloQPSTI06dk9CWAmZXXgxKEz/gzS2SsqKG7H5+OpDd863mB9PUudaEy9HaayG
MGSAI745NLd3Z8Cr+TD4Wo15jlIL9MUYgnCcFVBf/qmAYK9TayLveSBLcEjzMV0DI9lI65ijVb8m
eKf17aYbjXa7kr5iTG7qD+hUs6HGlFBZ6SXRB1c5FojBTcWksD4ldXfGHPBKITrRkzYuRE4IMu1s
Argw5kItgplyVCfgfMrOvdfIMIrF2DKNbOPzLZTf2X6hggWl38Q6028yxPYJsSJofHsgb0aIqHII
wEErK6WMwohhben5rPLEohXVLHiYqbqRBONhImcPpHvJ0kZLCwqwmcoiTL/v5XWwJK7VD7qTGLo5
nXMTCGQK7tspQdTzTIpA6b64Z+HlTIoir0NPqChDuXRhUKeRAyS10KnR7QGRFeyzdSldNgsA/M9d
dy7muaO5aoUZErM1SglsTMHPfqi3p/rCFqPn+VfnATU/O8UXfovCqhXzZtoEtS1Prw5dSs+YZ8wI
T6eysNXB5PqF5LsBz568B3uj8j9/U0Lh+pDCNVvJBqdZjH9O7pNlUNywAQE/4LmPAjNvYJGy1pX0
FpnU//Kifi77HlnYWlwE912o/HdHJi63xieV3/7KZpnt5I8/Z8q9vlrbiO3je25C/6Pss9pm4ITe
Nx9JHL+EaC4GtXTghF01fDHaAX4ZggwY51KivwkHsbZq9RLolKJ6K4NwPyMRyomLtQTqBuk/tniu
gV7QeTOfZGWaBU+4gQpwfLTRJ3IGLudnYvur7S1sz9QgVqPy4EktqZQw7C+sfsbWWdICLrcWK5Jv
V2WJFHDiD8DHjYw6DSRr8YTa1vX2Hd9gytsDv9VJRCQOHmT6IH6T9wimAtxeaii02Chcy4iPUlc9
8s52fu29asm5hGZcTUu8MqEfCuS4/O6gyLBSkz17SyPuxNvOrpr1J1vzTJoLMt6XvkR1DVQIlyr0
1KYjvlzIaTxzXjjJSahOr+jmJC2LPWaMoiMZo7XOKGccDc5Q4y/UOjhyWXE4nLTYh4zESvi1UYXY
qa0dcvTArUqgjkR4urt9Y3kcfB5r6sYURfo6lGm450ObM0OLrVNjHbGigJY3XeS8bRgRobxzAnBs
prNeoMGr7nxOmqpqLsvjfEwPBrZ5/okXbwgYB9d4jhSUFN9hnMcpFmhBJEAhMmACNr4nmzZQPAMs
SYuAE1xUIzh8ZJyetZ6Y9AQfnW94kszvZqjrUQy/MW+GIv0Tr0jzzlt9OGygfoAGPW2N8A7nVDFM
ny8QuXYOEGMPKzYS9vgfryfU6QFMA4sj2JGz6K6eORNrtaEJyX0Xg2gc+MXT7+aV4JE5lsXe8cX2
RTQb+bRAvzsUg0WiagUCKxXcMsSngOxheSl5wLmOejGTPaUimEil7v29OXPnFjQ1jg93yQbFj/Cr
40ueQHnQ0wtLlXL45aKsiTHBC2Hq2fht0uCCyJ4AVAbD6Lw9scx1KSBHOmuYdW9wxB4F7tW/WTRQ
DKsp89QCjY7uW6iR/lt5zZBx20xv2TMd1zHE/pAxWFiwpfBb5iNuMxUY7jHKQSv3qYr2VvKg110Z
T5lviqh2LTOq2BsY/fP/thhiPHT6TZtjGrDFy4TAubQvwsUaTtjRF+lmejtIz4aLXq38SuXvjRwn
WpJ8Bh71vAZmoSf4wHlBizCR+EW+u/D5WSqCr7hqsnzITQUSbBqqZj2USoXsAzTcAdkw/mQu0wQU
Tna26lvQJd6Lbst+HuoiBJbwiFRrKhfpoTKjjRvHmSKoq0MVrzRvm2kvT56G2gujbU3gxkFQjE3F
bpVXCiG3Gg5NTYy7/VLZQ1kIJJRWt4Ij96P3UHh6l9O383QADB1YOSuScn0pXh3pJOqxZXAGzTWo
ACv+GdEjJKwnGLS9SU+S9kW3G8uihkuLi0Clr2EgvEuCIcmqRgdg+rFuI9gAglgq/O0yiujozZDj
nY73phX1kbRPIXVMZVr4y6+kH92jsuYQjIAj21UhPUAzO7Amp4mGtrp23NG9auoNSr8UrrUTqMDH
J2z3279tgpiFvlHAxhrRdipy/RhRRpLuuWp259V1bRI9C47lzpV4IVkoRG+xKFJCob0rB2E/LKNb
Q6VUtHBDrT6xN16k69kGx3EcVJMZsuQSyiDiIBb683Oy432t+RLftFRff74At6Xjue89RE+glTbb
ODavWY4LNpxYSavJhIjFz2CPbbVBBlygWkwohy9BqaT56j1IlojPPXcDKzsKuJWyFDk2k2cOjG9q
jCLaxAvRKP3uJ2139brt3tdm/pkU5Dtd4rNMvSKfPvtkSwQ/iBGrdMg/X/D1wBd6q9FaQi6d0y+Y
cuPehkxP7Sxzs0L9hn1qNfvCXJTGlSGdZyZn9tU7DJyUvLOBvIq22/qZVLqlwb9wvaRUu24LsBKo
/lzZf1WugxxkWzTyKpQKTuFOCSW5ikGCDVxn8Qs5k+nf67hypbP+rQKQi3WdoQAJRhVPwxA88T2w
CTUbaRBiMoO7UL3WVUrSAza28zGgFzIxJZBKJgu4Yz03cciBR3UkOBUp1vrRSz1juVDeOpHMLcKm
nG8bCfTTq7Ke3C08oDaWBz0j+3NZB4C/nPB4gaiIZgoFoQYP6ilcvNjDUQLrEgzHdkP47TQdiWyk
TlIo3LpafdznMa0IA7U68arPOBZLdnniacc2B7YVMmTRD/GYJZu2P+j2hpnzWFHkkphcQWFhKrlY
B9Le+VgiIM+xM3fPVId2qKOjneZL4F+tY1zD5+/EfGZa9fQaMKMiYlXGqsKoL4Uv0DBMEi/8gotw
CXhRYCNiO1NZB2C2WZW6gre/xyVCVBT16LTC6yyA8uiB7BEcnHugYIS0Q8DzvyaDizXMFtR47PDU
JoNgzIZxvv0AU3VZwSBFn2uE5K/yJN1X4Ps/4Cz5HsLfgCa4tvXAXNtQrSjioGDh/aHsbghZd8Uw
6g73k0rn5Mftp4Hfm07attm5a19bX1LpF9fDoPoP7VITvYnspbHNODM89IdN8lWNSFnIKb9vhxoR
4Xj5t4iIuKSCe1dFMAEeBm9TrQO7UNXWmGDl7cmn6kR/6S8ew8zM/oyY8TsVa2RxVfRxtYEZCfW+
VeVOkpJBT+nc5hEOPJuCHP3yRCd8STSUdYHnpIDVQraO+5ymDrp10xH4NTknqqC/C78n7gE6Fjl2
NXdNjfe4mUmoeUGpv+QzFk1ICD2yByWStY3P2Wona22q67dlTRUQYoqi2GMlNoX98c68LuUY7rXI
own4z9xgcFcljhDXBG6vBDsMs5IZ8Uc3YV9oX0LI9LApLda6sAYqiSYPAvEmeCiXsZH7LO+mFIv8
5QF0FUu2Bh3Fa9uXq4/4pzPKNDqPBiLSdXQRNzVzCC2tRI5qcWwQyhQUYtJrvy3hNt38ARzbSEmF
MWwjfJDpdl3k6RdAqz6DA7gsfxxRw0S2vzgaKMOMMo4RLlY2HEXRaMhK8kpmWcaeR6SWHHt15LMt
lRV01wVexQnJpHifBvwm8G7ZbaAcCiMV/MK6CfuDocYD6oBqG8FHdmRqX3zg4Cg9w/8Bw3xEnUKs
QHKz45UoFX5PKHmoZK9m6JYyjEBy+L12oyA73XRAze8vO5g5mKcut8USW032NBAFJQYAQBhVHx0w
4UUlwEUPjFPmbItlAvA1zSLurcmWYTuncSHoYheHX5dragbY6vlox1bfMC+DYdx1JigRlj9HPctw
rvfyDwGmtMb8ZU8jV2dIJx3vWVY+vWUy+TmZpfZa0ZV8rKuIDANZZNShkiCsUdDvjGJ12nJWeVrs
r+VbwP0fA1IMz+T3H7cANJ9FG362q0mCt6ZzCobL8HuYsWaH3JtB4+IBYlPzeQxYzANV/Tto9Mq/
DdKnx62dC4xJ6IaKKyclpAcAS9pCAR4wdu9o7FecJvT4n+HhOWQZkH9myWJxK774tLg2WCdYLpio
xoj/n+dLKYXNTO8KpvWNUDL9XOsoKjvlJvEDF0b0juE9Xhe/F9cLSwY+2cERlGyfJ/UO1Tl3VTc+
YLZD9LQpSVP4DtLRcoBI25UpDJyR5/JC8dS78yHM0ffEI3mJHVqbQ2nBK4ZC62LwYCOgkz3tuzfY
NXgJkPU/ydvGjRLZxCHjeDcwwQwg3wZdTZZHofEPOhGbtxR3fYculxhrbFZzn0d7R712VhKNkLX5
Q4y8dyNIMSN+ZUrSFTf+9mNWI+PoPfidts49uq5FiLdDtaBz5QOyXcNz/x6E9B+4SaEr92inx4R6
nuLW2RKuFddl8PyWT//nIY+P6fySwcVFsDQMj3NokGqS0dXcaaC3u8saB1qh51NsmsYZPBbVrqKz
uNiQk8M++91prIIQqB8J+ESeP7W4xEkdGgWdcQErsgUyTuU+tIIwCv/YlxL5L51kt/+JqbuBAk2w
8cITQ+LE5Lrv6+T1s00LjMPplDVYbvpcFJFbgWDXYzuEdyx1fciQNnFRlhlBrimdqEfW4ffJQviJ
bDSeTFM0o4BpKE4JvvyuYaJgWJMqIuzkDLk9dRNvvNzN6spW46ipbvOG6z7djloEb233zTTLUQ6L
f8bxj9Crxyxb8DuzCpOml/5VKJBhGlVPP3Bwe4j4JTRPn2aVMVbXk/9KG+06Dphc8fxtV6wHvUWF
Tl2MKJMLrs9+z/49QhlaG6w2c9ZsivSoS/YW2mdVzJfWBTomgOX4XpTWKSGSlejG9rSFzqJVH26v
9YuiF4loRgY7fbnbtQodOEHbyewMbytQjEt0eOPEzfjxV2aX3R9iCiof+XeqZ+pPcLh7QFVY11Oj
IFMnyzMECXJC2YSdVfqvGP8OWqSbGkzGnP5fPS486bvi28N6VkiUXIkP7F2bP4Vafn02oOLJ20JA
X9z9F4nIoAeU5UiQH0ab3/uRewbNhp/ak8dG3nXrx9js36vlDFshiuNedLtdZGBl8x77N/C256pS
d0rM5dzyMtvFzT0KgmiIqpCY/HxC1zO4TC7OnVFhIMzS8dbwSpnnzDs4Q/NpkoIon5mziUiU+ezD
pGdQnc2STOSU6PbjJa0uwBo4EWHyWt98X/NBc7WQ1GqXEweVNiucx5kD+B5KVphu7XLDrNF9N4q7
cmTIkmd7PwvYXM8cv2RzPorzePfT3rKBM32zG4vcMOJlwoDKoNJCDIZf4wtbm0MeRlHsn3iDnukh
9jT9daUEZNLVI1GqbxNFR8itFU+JcQyJul0lDVd7NSqu9NAKSlmYvWszLNrscLarbje6EghL1PZf
B7xwe964RmvD7RdXXwrzcmxmoErGU2pYooCcmq6Pn9t3CQ380vNfuHNlje5cXh6vwOkhYwtUW1nn
P7y+dk5VfFgoBz5NyP/qTZVnjQ7O+CRlviE7qcMs13hWRHALLOXy/oJ70Lg1Jp7QZpv+JAkBDiOD
qzeHeE9WuHo1hVEche6iCLODfGrccSHztINdx7qLPYDiJyJWSu5Riuac7CQggXDfqYg9XEZZo2ym
8MvPhfJZYrsSMNcIERYL6RF8Ps63teCaZJus5UhZbFZTystiTUvle0q1AVcZjvAPzaUCqz/K7wE+
EVh3/BDPxPGgsed8tqDL7LO9ibxYkMlFSk98wdcOcnxTxSXM3QOVSQWWLNccgBDtvUi0JS0z/h81
IYIvUUcQwEH7ki2wD8sGrM1gGcby/LoLJWDYZXmalqgyP1frcwrNhxBFsx/zvuMCzNsQxLuol7M6
kM3lkt2k2FiCvy2zWePzkQrObiHmv2B3VNPiHBxVVqWuRdLfPUs69mcjj2WvSecs+PLRIHXOSS5j
HUowO4JR3Tgrtzjevsfmk55MUNp1JIZaOv7nfJvtldFjKhz6YKl639SzJZugjlk1900n8zypNTx0
rbR8ypVkOzScrvuBafjmAdb6BH8gT32Bb3GQ4IC65LymuEOxYFjWtFECIT6GSL+vS0cWvLotnfTf
f6vTqzxbqJ7Wh+jrwy0AWLfDtFbnb6fnY4tnRQnvljEk0avVgcgTJQC9iPzHqniVeRh7tUULVCPR
v4Mvukl/Fc0AmFr238hxhK9wAHVrASkC+mU0J4Rlx5LsM3CUv1Biql26K1ZSX0IxUcOTfEkV+EMx
NXeYnIQAuXD0Wt+SpJztPeg/4akkadSzFTXehYpeXD03xhcWvJPwdbJio3ZKaaN1Q0tIWHG8BbX6
kHCUYCaoBwDMASUPg69zfXKGZo1egXJUrBCWsC4vJExoRgLIHAn7GFaNf/k1iQiARKF9oZpQAIyJ
5F18aVKit8ew3NCVk3KdYnTL4ZRrBhFRdHN4iPIaVz6rGl8rkim222wteGSTP41tQec4sYkdVCEf
nQlph8bPhcowY0T5ftMgLGosnl2Av2N1FRqetxw4Xuw/EJqCS4UAlW9wlSwFcdYMS7us6TasBBm0
8i1HXk4TZ9PGcfB0xDQwoowWZumdwObBaTQW3VxW4ogFVcm6z6lBmJoXdWdszXY3FzSorFr+tDtR
dHXlZ0sUneN0CWw8029c4fIKzj4n3mz2Kh7eBc+2ebzvIb6w9iv5SuAD8rBXUF9gdslwKeckkP8s
JejGK4hnQWuLWIxDonb6b5H2R86fJaJO38P8iXk0eBe8av1HuPEW5Y5SESMgKrJGM9a03OI6ejnR
2lI5eaNDlreCTI3N/Jfq3Wc/kZKugI0yYanMs0q3xM/jUCDb5IvaHHU/HeK3tRaTi7wUrvPeXlGu
o2bzje42ObkTORb6/CwnfQ4fyLcbTJ4dcrCB228S4k4vs4HFkMMZcAtEbcBcEDyDq3RNtBwhfefU
R1D2v81HSrFQUCgsvUj0+X7CNpJvRMio5izhEOqFt3nZZbxmz7+EZNnLX2baLo+pqY5N99NFGP1N
Zm7Vnfwa4RYhsY44y2bzsOaRYBh0IctK//7F+2Az3JArBuuWMPGdCE+VjRBXGEyGQFR71sqJQTue
YcGCRk/TK0pithUEMe/iNs7669m/rgyH8H+oSapBC3lTy0c1DjGFKcNgpGxlWY/mo8TmmzEyBhjr
wRoCMujv5Ry4B8YrMauVJ0x3sHz86hKc0H+s45OfUIMvetJRRTUauTu5Nz7Vft3PeCgLZcDRTeJr
o9avuU4UhEQ8WK6A3Iw1aHbbaHTGEUzuPvYDRF0W10eIAoqNgnIJ4AMjrOr7p8MDEqxtyvBYbmrG
N3HpRVEiiM2K07ARweywJSDWeRFrCCVJpiOGqrsw2jiKrUTeWinxPgwvBRgMVFkCGSbC+W+vbFQE
W6zkQQ4HvfVekfTM0nul9dDQ1aKAU5Emj1V5MNwWWztkYxYTlYipk9+M1z2wOSBxf9bgcGv1gJKF
WgX0LeSFy16pBGdypHjVI/Wv3Y/XeQsyNL5EkBEoDsO3bzwTOgf2rFmR52u5MrsFXmLGzNt6yOUZ
BcTsBtaBkS2hJYSSSakeVJhJDnfX7HwtcES1x4K4pj+1ZjdVZd6Gv2Xw7xCEbEgwvWVCoEKeG47K
zW5nqSSdtLHyV/rBbMNz9+Jy/n1FTLnwhP49IuWsXD8bdPuhTgevUMWfT+/3TAHmg6b+VGzFUrzV
bbdHvRJrYEanyVR1xwpAZC4ndNJ2L+X38Ny+psJvKR6IVHZgbgYwsc4aXMkPUoRZXLiJZK/LlY1E
Li2/TIjlvUv1QcfFdAzAsqHVvjtgRybqCpNH7wfTr8UE2n77d+luAQ2m5kEl6XrxK3f7ngubf1GI
IKPzZcyt9odL6g7dTt4233WgHpvQFsBYVMbEbt7bQNZK3/b/QOPXVIEpnt7zekmkeBRmsgX+1ZtA
J4aMOKYZ58gYOuoY/guquXvZ1P5aRJiMeYeZAiYhaPqXivJ44er4aXgXzhhLNCiMlC+ITKni/Zyr
8YXHbFOPshdo3gqZCDqupvCCYDIsT0kHvafMyripoGGoniBk9oTscP+0Qg0ILY5I0ElqlBobdhoM
8RNQHNBiNGU23rGRPO+TBnmqzRnOlzXKWVjdDMnEZJ3/kN4jZ8kGVM8Jfa4ODrb1T9BbcoRMFLaE
l/PMZDT0ePeC3rQYITPztZUi5v0R9UjqiOwfiw/7W6MHek7j3htZIgtPJ+WtY1TM6JEzCiNATwhL
7BBP8EckinTW5DpXA6S/tIHVHigbEAY192J3BWkZFnBp4ECXkPQmpW6sfoOmV/vy0GWG+HqlCz/t
MVkhbTST5SSYxpmGZ3Xe1GgoYx8ZsUcf+n+mf5txgAXXUxr5orw2YAlzbTDzdMiQT2m9f34mo2DF
9ZndK+QVXL4u3I29vgXx7bARC0Wv4Ly6qUogIz03PP6LbKMrcrvoFquLryQXZ7oNrjXes6X8MO6w
JNfmpDzYaY3SKHWLL0sN3fanuhtPuI2Ixkrr6RGGLp5fFzNMMcd0g/33u/pLJjB0AQMaGVGM4dCc
lIchL2DNB89YBVc0Qk0/cKllgGLlV4XiuY21tdyWWxKTkFE7PEYwS/Jty9H0MjcA8hOdETqJxMdP
IOh+xKeJXQWOfGvUFr8xl34kUrNklCZQSskbw6flnVOHWbTzlKqTkaRQSUYoeeGv5qnM6LIx9S8n
nRSqorwvwuriqg2srKFMPE/crgxMr0W2AABzKK4WvJlIieMbTS0z8u2/Lez09f4hFMD4JpJGl9Mq
sA2y744VOG2HEFpl8u0AlPaXzcRMKSZq3VLko/fALk3kYAQS1U1eUrhzxMueXRAi1brVpck5l/cQ
PCfhfNdxs6GAXTYI/G/na1OB9X9ZC9o3gEOiuNebQLXwnnTDtMrTMpogoFh0MFw5M0to7kCe10aI
HMS+mae5CgvodccK0c83XN7a0PaFF0FwxDjAOkTCz+zIAqFChozf0rL816uZyiI+PEV7dsrBYA/C
lHv0AxZc1wcurBVrzOyw10B8Cu4ios+9RTgosy78OxbfEvgGpVoFPaSCbrhjdtnbhZsME/Em5DQZ
hmb8quJmC8xd7XGe7n0JjWWAAZobm5ibRnv6Y1yTIybn0+xDpRQtuLpokGmcInXjhbZZ3MklZoV1
+rpJisM+T0rc9QvrHCtik+oTfS3qoW23lF8KLwjfQ/ECFGDZ10gLoGO9PzmBhicxgDsBfJsxWzVb
nW9/aUQHCAqlZeqyZEqKhls3rUvtumaarYkcVyW7VuA7yEYJkTb4g0QLkgZ4EdJ4ZVTw7gSQcWGt
NhqIbAiqX7i3YOMfhJUiIOrA6XHoeWK1aaqzNlWSN4S2s6l4qNUuoQTSPQ62NQqpxHoo4TlZIwhv
4xsigQAMGBUaEnnWRgJvH0MstkXZBlug3ba3iiE1QN1DFMSSXsZDT9+47CGL33PVWDc13QNLEr5h
5FYph0OSUoBYOsf7GaOjSgOac2BsOqy7+RjYOHO7NmnM2bXWkupRIq+vNN09ysEKmgE9WXRAfbFa
yFlybBitxepa8Oc6ftfRAD44NU2+OPKKi5HqYHyTT3rIKpu/NjtlUAturb7PgzQvWvEIM++NVHrj
QA28zsfrc7SMBdR+w3mjSvn3NywB46HbSFI8Z0/RPrpeETzuglIdbCXo/g9ljRXxpdNe5SAQywwY
htwj9Ux0mvcqfvszDcnYp/AKtPEEuk+qjzZY9FP4M7IOCL/lFJpFLr5Dg4L0zCCOnwhEoeynIOUa
d9gilxY2+qUdri49yiTXMYQccu1kj2q4KEKGMspjj76+SEqDyZ5fSZV/jWo0ROvM9FqJ6nQ2IoI+
AyUMaYAY3rvhFoOvBG9GqdxltwPIWPnP4WKHpepg9uAzx5JRlTjlt/yT1Jsdns0KRooH3RgCLJtA
UhA4Ta/KtR/9y+1DpJXvEguIntqfT+NRWbImAOsVE2nSR+D/kWujYSEs/wCDWE6cQ8QBHRhB6omh
JwY4lmTnp7cjVPNtdESpyDsn2V9PD4quhcYoBzGFuhYmD3riSfYTyu1SYvLVHBf4ystimDXG+DAL
BcrpVvSl5NUam//IoSs7MtuF3X5Y8ifXy6pNlnncnLkYYmYt7AoOBKQi8Jm0EXdMH2sfEQfCg0ba
lIOlqQELrq6qB/g0VVOXy3KxUpIrKfSZIXSTnqnbyUAYcNSgFZBh6VW0YDSPpBHP0GOTXrK4prjg
4ABXawsZP+xYr33kAnfE4JjYWlxjVgb/DOInQp17Euh9Q9r/Grnq+oFSx/FiZzaBtIAz+EzdCRkH
w5o57q5Cc1sWLgqvKywEcbNbLnrw43aJTpalS//+6Vz5lgiln4H4TRlxzix6nZTW9qWFE8CZZ+hm
MuaYrDshZfo+dnA87B3xgIV4uSShep0YaNVu6/6w62axA+PLV+TaqCTjcEwkApxnFL6WmRsP5fsv
o0WwZiZU3N+V++A77J+f/1WcGNYPJJyH0ylQwFshF4H0Tk56TFvBnqDbq+5oLr9jKd5cXfdowGhK
I5aU5l/DJYMnHBAPYp9tFRqb1qckPNwo0SNio45v1sDRuvYE01SS6QlO3Vca36vxSvX5Yn/2p54S
bki+E8L4wAGOSDb0+3PaKVxuAynhY+U0oukJVDlpAPdEj5Csu0pKOiKgUdk+YV/dDANhsBEpDEk+
XvSMVsh8NAKbH2a+HFaBB8Rwu6GkA/DV47ePdXWqmvwckoe9FWd8HLqfbHb+EsEN3W7vJ+9RmQNM
XRPIORS1aGssic9a6bdJys1nVKEv2sf6lqITLb3b3KU8EcrUoTlPguB0qI+vnn0Rq8HA5X8MVKlo
qGrc6zdMDW8KywkySctYsKhh0iw8UwalWLdn8cwpkyqO4syQEVtT6n+ZFWN5DGqcuMxW5NR8aNTi
+26Caho5QknzsSyw4+ehMk/IFY8nrqh4ew4r17y78uCE1C/b7++B2T3sOY+IgKT3Z31gZopHk6Qe
k9z/CmI/tQ4+Q8okTr/tAyZIbwkCc83ZCdd//ozUFnwZGwF5eAlLfv0N/hYGCtx8MkelaATuFM70
lBXmUbhuJOiY3JdyVHBhGGjz1UUk/Ayp8aFgqE+rZfycSfkOv5xcA4c6ECosG14UgIJTc9Tdni2Y
EgGoDQoKcFBDPycTQSokaIZAr/Sx9hLs+3i3lb8RN69oq0hyasPv5Fr7OBA+msFmUog/POanMEqe
IJGU436u727FyaL0omH2t5u/U8jCYoTpGH5SLDhiWomcrkFF5nkM4hExJ12RatkXbYmtLJaOdsCb
gS1hRMOvnNN1X+3Ccgepz7K+tv2LLuQ52nOdg0+DKTcxq0VqMGb7Uc1Ep9c99iK5uwNXAK9S2Kwi
6ItQ8yEa8atF1LKs1WOIxbm7BWrwHQxa7glC+4vRXdcHVqAcH2XDcYUvFt6B8oaVWeffrPWZLkGW
+5g9nYhVujwnoRISyFoorTU3gm7aTwTP2CEH0qTiZHC6mNnxIhfCDW/BGvI3MiojosCQu6epmtzk
hFo4Bos9GYIWrSvMnfxuJE005vAUr7E/VrdLd683pd96F7z4AhplLXqXRdDx7SN5t0HKfhmetV0h
oln2VgAOBkk/aphJNVeBSXy+iJFkfAtAbDqmpcKrSX4sbrgsTFn2Aoa4KiJp27ruFtRo+cWgZu4p
sIi+VRBPosUPyRKxA2FVH8PlMv8iJpOG+Qo9O0r1i7xhcNh3pPsswrGjz9iNvgly2TqTBGkUKrHd
p6mh2O3eQaX5J+3ZO0Ze7IAcu60ENE32Mgl5WC+7NB3vpA3Bh34L/MmvM+lBPfyEDLes88zm7Has
+ajkG1codMli8DxhrDDaqE/7m4/8Ulo3Lg9pGzQBmOSv/HBS/WMFfIT6qC3mj4vtbXkIKH42WiS9
zsTSnUgT1tfnEgBtgMfk8WSU+MmOa32myA9HCtKi/+Xh4uUamMrLOh4JzkKPUNshcrM/155PiQXX
JjX8SgQGDUDOuoT8YL2iaWixRhOSQmd46GHe+mX6skq9bGmr/GmAuhmwzIOb/OJ0+N8GzZmu6pDq
m1oQrMMno826I7BYoZvDIT5zT78UnJTrRDcGNR4xkApoAXkmW/477jttv45Q6+FrYD/8dfk3sl/n
kM0/ly8uKoWT1H7i7cK5+4O6won2yfjYmQIntWFl2wPFlxAIV5b8SgQj3LPYTJ8eHPltjdfWjynK
SXamR7mhcD73CYbcil878XwOWNOSQocebwAutnYTeeBpS+pULXNVyfB/80qjino4qTRGaLPuydh5
0CRSdRZUAAz6lIGD0z9LyGWHGBjufk8GJtcUa03on2Fz04WertrJ8PD71aDtPAw8PRohdcQwDpAk
vTgGrUTEvbPEWNYKmLhci/tLmBkm/0X/2fQUNHGJ8FlQxRYFhB/d1qEtuXUbc+NtbsU46pYkOB31
/IPaX0mAsKLSPn2tMqx3QpIun8qj5aD84ceRUTbSGGoVZkFvAl73WhSKB4XIaYGweIsSgJOswyXg
PJA1mk3/GFs5fZQ7QyHaZgjLlHJCFxb/8EXyEGx8R86v71ga4Da8nP/E/yyzrw48/cRCdazl4hLT
+OvT4Ar6OZFeylsM09ZdSI0fzFLI++2ekqclwMdBUkqzlt+YOWEwk46pzqcPVLonpYxVIRjIDmRH
bxLdnlsIwjAjOVlhIcs2L5CTwJr8XBysU3EPZb2d7/cl26l/3G8jbsyQjd521OWRbpoLHhXPq0Ss
43IkL5e25vPSVchQbtpsztCyzOrnQybucLuTXj4N0gL4mof8WcNfzcrj5zB4gLSXhNTEJSQQW2v9
wOio1AaRJOfY2+W1l+1Tf6VdLVMSDVoSk6C24E/1dJoGo1l/HM9VflQ0uyQVcORLpZWH/b0rW0v3
NhkX+i2XYosq+NXU0VftS84WJ4x5ttAOgaOAD2zc1kb8rIXpWYTp9lXAlhKIA/ZHjEXzIMsTRPYT
TKj1QEsIaS4AasHEi7JhNYE0jHVzU+mCqBKnsW0Uem8xe5OkJQoJvGdgJ3Mu8u8IAyM1aPfw6P2m
YyPFKNz46Sbcs0Ny8/vqZVxXtqCHZNltjqJyJPkvtSEOVqXnXWf1gGFdrl0ZWFtsQFlEgiNblizj
4BoSA/BQNAt1ScApFVteZ2iBGKoDVXfIYYPt9waw7NqokcRSzf/gov1CEPaw7XGFJB+jjFjgMgGk
VK5R8kznlVVrd+TB0trw1pQ3hmJ9mqGt232jvcwQjWAec7F5VaOzL4wPO2D59KRZWDa8ggVaqb3C
C54aGw07VAUrO7Sw5+Rlzc0kzZ1b9IF/15VX/BTB3fWxZxvikLiQ1G+mQEjlpThcLN6U0bTRuqK1
6KfktaOBRIdPaIyPDhQ8zN7oDo4TaWGrACdBRY3OvheHM2fjgI7Tg+N5gUw5UjKU23OvbhNvn5Dc
nMyuZ7Z5heS1T8irvSWtcJdandxL+a+NY/4O+m49deSElTJjUESIOTqrygSRzdtT4rKV04Bhfdlt
Iu52m4g++zXAfZrDKsnZwleSf4Ze47FFHFZWrHGUup29Fs/VTx0rREqJ976wxnJY+a7hYDNvBYj1
q/9aksI53mI/hBOiv/ChwkIwSkiWE7+LaNX2+xxggc+kQrGFYpUmLKc/+iirEfxYv1ZK3RurCZdJ
kPWJzz3c11Y1u/WcqcTPWfA04VEaiBhy89DGnyYUoocO8s9qGkMfqJ7CiwlvdyJnVh07LWG2TkKO
qestlyxBYa18krNU6Hy9Rpm6FIt5y5JUmj+DiSfNY6N/eipG7IAxrAQ3W5BCdSyDo7babDJYgGZM
4eNlN7ZZlXQrqip/F/6XsMMRjkZkgF/Ogt2YLbk1jLvsBBkPNWisSEdCb7CyHvUuk7yaKCgLbay3
qWLpVyQhVuG3d9wTdxPWJMXPiXnP+DKHMnGrdjtRfOp3TREIM8SP6JwN7pkimUr6r+uTMvRLl2WC
HpvIIWcvzSSjsmBdQS4rcIJw1WNgOC+RHNtHMBMFYi+1O5QPC4Ipa9TciZ0kXyFdCp/bozr/Im/U
M98LtcnHWiPdSe1wbUGpWrhkri5skEtamFA8us3c/3EJ9ZKOHzmd76Bc5vk8HqAQqnnqzp0s8kpw
SIy/8nxzTfUrdZYSMnYTOkbfofPzIJmoW4fqnwqBBtkL62/zHYogHrq5FdwQdpFvpEF1k+0Nuo8q
1eFzzwOA/y4n+tDQm7Xsorgk+iAuUH+j/obuefqEPuPw0YrDKTVH3/acRehgxmuxjw87UlUahAaI
PW4S9Co8jvXUUwK2TECsFXA9lP3OwrIGCjPH0qtu1B2WUzDPeJF1TQrvD+B732FFgUhaOayo2QY7
nFAY14jTaP5ry1v7vBJIIXX+05YH2xnnW1IlvLb5cS01nyMGK9ozX+Q4eYJ0X6z/jjKxp6R8NbS6
1/d/mA8sjsMOYDLdTO7yZP9IeEw1EsXCQ/UD7XvAE5igKcQy3zQoSPiW1PBvsDvUPVPDscavg0wP
ZCUDSdBr5E6pqxLR8e4Vtatx+o3nLaMwhhqQCZOQDWeB5YJ03fQTF9ufkYTsn5T4xjlAzxl3LSPe
0l0Ub0hvdTWxKl0VLmo/Bewk+WQ7YKilIB0oFsGnYhPNMyEa+Tcf/zgp2fQM09gXTGcgxRB/qG/z
u5W/jrOSxiK5dgikLFV8fjSloONOhcHMgOx8QUtycO/PYY83oIWgnueN1lposu42qkDkJLf5va+u
hsCrT1IOQadLFcxCkQp9yOwjfCX9sSWiPIuFrj6vvDVpt6xPm3FoFrsA+1bMAG+3NlIiT0C+8bd7
o3/3CmS9CiOjWTIWKOeqlWfMWCFKD+7c25uR497PNMO7q+uNb2llctZvdXk1CeTkpKTNjKp2/kJG
QghTIqLR5EBBiXnGN8KbkR+VErDeWI0tzPzCEtZ8Jgh7Bb1jDMeDPlLbVZuQ7sZeyNmwAC194DgU
zqRT0RdOt4//XAC8EL+cJh9OU1at6d+Bx2tL4QWR+xtYD+74KvLn4r5zVHypT0Z60AWri0U9Aalu
Z757V61K0LIJM7BcM3w5fUbbZSOrY6ZTcz43+2EnNTVvC/USPRuVAS0n+rXh8auLVuodqKg3B0f/
atKnbhX7MZ1Nt9KdJ/LAPL3ZRNtkJSlOIyVE8dg/opQ/sXt9WUbYFQOYdwPxAIrwaEb2W2AUf3/X
0g/7hMV8pqyRQNNuXTbeWSchIs4YN+VsGWQMh6Le1wJdsH/mq7m/GHA0BqUfkCxoXhBu57R1RD24
8xkXS3+dq0Y6ZRG6clyRF5Ba85zFRkFim73PNYg9xj7pAKU8sX1EfXJPpj/yOkPpZ0AwQ8LQE+MH
rJIYcHTFsPUDOtucdVpKIN7b8plHUfXR6PnSzPXDuxFEohIqbhMgQ1gLo8EaEwl9+Uax1G2pxw+W
HsXQfQA8A8OhQewvSfJ9hWslX/o52vgaoJbFrqIyo+9Fd6qLjyOBF2mrRMxouF5CHMJcbCNcFMZQ
2mrsYWKTYqcj3IUijv8w3936k3zVXTPn8RkJTftbiX5Ycgtb65JAMAR5NrWZp3kYRwNmMRQU7+Ha
gBzm1p6cRo0ra+dTugUPzRFYG6tspmlOgIfArsEZgQKkWa9/u+Lg143yJ6ChQy5tlByEDjU54ytu
yIv8sv9nED1gSr7vphhEUrpEvnmBWWpTX2YuyJ9vnTIz1JHhT8bBK2YREe9Jo+MTNyQgaMEuqneT
vIKkVtcue33VQ3xRAGBBmiyxXc/lSYE/wezXh3Rw9Wxc17+QzEkm8he8B4LWrpDgptMddLtHHhy5
3qws/BxOipeYHXxKeF5Vc8cWdWo6JPeZdlvF6wa/0rwN6i0e79dgWv9xF05tWmdoOYJ/e/K3yzeT
4TF441W9pBIqz8uRSUYsQswqOp/LpyQz8N3TNN2yyE5C5g85jeHFU+SikFsdPKePMd6bMwsyYR3i
XaBIdUTfGIgOdydXD7ut7g51QowyrWZeQqW3Ih1v3g7duoJIN7ZeWU9iIWsaI5PR6614+iTiAmLG
cbPl7ObMqwPAlxsHU+LqqcV/opy+a/nBD1JC6bPf3H2kj1gmXdn0sH91Jw6oaouXM3qA3JkmTTRg
fQT6uh+/Y0kxoqZYyowIL2eXSQdwutMHIj93c1AphAoSLUZxm3/+YO8AyjdWZc7KhYbaJlUdFGwM
a9ofMj96ngZuH4T+cVcVFR+R5UE+GzGZY7/fYRlRolvaOZv68+zlcWHrNjk+9oeLlz94s9/XRRQX
i0wUqz22rkC+3CVs1bbd5z25QkPKaaAHMwFvhEZUmOhjFq6swU4MldcBfP9ARRrybhWABJgKa5v0
XslZaJwyjGOpZ/VAadOE0WoB7+AmN5QweMQ+1TmBGCM6EBAkWtkmGRdMtviIMUZyJe5eNwdwYKqa
1PhqFVDq/C9i/9C97u4TWh/Zsh7R/6jcOM3CagzRrAHBY3AvyS097qZqz+rfcVLnYIYCZiYTIiLU
0VGEaJPIkGYdMbpv6g3q8nNL8J2gh2y2AW3NBk++rYdqYCuH+FUXFeZqZOSY/yXRy/nnB87y3IVY
Do7eQf3UbaAabniRhKxI6w3kU/LaDVpw5P/Lz8cDdG6s7gvwxBLUlf+q/YPeJVtVVMd3mmyrzGQJ
cvI6I1eWvEE5X74oAnSakuguc5WYGQ4oJoV9vk2xYqkFoLnUU4IS/s2/pHuiLHFepSC0M0bWC3DP
SWC2Iajx0HkHEbqFAFbRf7FIIE3NNSIHBaCsmtJTBQPsSfV5H6cPinJ0u/tls2hMZMHVvYMAS/+q
17yynuM5SeJgdyTCT08NXkz/hWWuGiQoI0ghc0ww55c9o2kc5n4Z6KI7OF/Ax6faj6QNHwScrQEf
AE1IcqmEr1Rf+z5Uokkd+0aA/ZQj22ma56mpjKd+bP7nLLyn3RFcJyVTjzIFsksyF6qjLrTfg0H9
4uTlsl02/mRIv0uq4Qf50xnJ87HaTR8JDKCDivyejQRRYWF4sRVW3JylO74efFX1wjo3HCkhXJXR
9kklqPWESgZH2SfRS7eKWd0bI5cP4GXHAORQjijSPP4VsaHdLxFw38X1mpz/PmaDR0yBN2hdTM6S
uc75UKHI1ov96M0oNYioCDVnWkDbGiAUX2OhIfMUcbDuKNkOlU5RJmwoApPfVwFHPTMAn1FIPXuq
raIh2dHczmujQKAhSPKF0Alg58YThS4lpfh8rVvA1r52+2EaoXYTl2GAqLT1C95RcqmRW1eXw7Kx
zhVpTSj/JbLKR53/DTbXAJhHT+UoCmBuPlTv+HcrktYfS8hsuvkHyZ+4xmPowATwjjcMYIXi/Rwr
PAqc/ANknBX25CWH8cxzeQy1ke4Cy0FZQWzPt3WaxS+eAtU3JbLP9QO55FtjqjrjwcPxYPD1Lpaq
R9X1tml/1Ve5sQwNTB1f91c3mcoy5dtaIQq/PafAcl3AfGCMM/Q7r7BQblP4hJMVlxPOh9ekgiPO
OhRo15KFIHog75HbZgjLSELvbvXljK5PXDiqlSwBDt+UoWy960Eiq8QbHyR8tiTk37fzEhLjndcl
Y6JEuiLLZHG3WYICQw+Lqet5tuoK67BdnbG/fpH3eYgIHj0v2vPsMwNQSVIoRWvIZigXcXF2kGQv
Rvus40Z6qXlZCmV4gel8l9YZoKzdUFg8UaBhKsUrbm6oJtH/agcwpCM9CC1BA0iw/Q2V2zoXKJef
hH4mrCYWo9TGr6zS+UTkKOaEwMvEhMktUh3ZQjgfkBRV/wqzmexoKMmGv9I445lXjUHfYFwsB3XB
+QnXdNtMoNw1mFZXpooKEhxF28dcXKTok/DpKbz2lr/gSPEFyu/XUM1WcrAM5e4D69O3TbHqwxvv
prA+t5fxDkD05th38CosWK1J7VvQoS3XJRa0+05WnTjsKvD+ViBIK6rvLB8098cOyVRdLl+bXgAs
rCS6MHDc/uRQXPfYDUDg11rYF6JJ0fVWCmCEjnONdgV4et9RyHoKtLuxfaTooGaZhL3btAjvuObt
35I2Dk2AMorHHgsmL8uUOdc9MWgQkeh+XU3izHLQCumYj6rU5Ii8LZNEPwWu32Zx1OJRZLYZ4GNX
UgZoitbJNqMcMh0ulF+Jf6xFMnePyps9ku1Vyose6HycSWfSAMrU0psrtGG8ZdqZHObMkr0L+M1V
ZbnYSIIgtzFgvFMN+qxTqs+gf9ww8MnoVsBOR/zz7G8Ua6h06imkSoWZG79em/7bB809oEFTsArD
WQr0xPxlCmEOJR8gJgwKXOzkDetT0nUsDtRHFClSRGE+FB8AXuoFj1IMB+x/crHOagEyi0dT2ndj
Uwb62POVS3wk/vKsEvdDemBPJOrz7CDWhwjc/PuIazkrmawh7+7/CDlGv7pRYlCMec9/PQynmMR8
L3QYFZtxbrep4RBmMuBZicS9NSVkTQW0B+9OYqxvI0jiHh6BjcEpA7titfL/bW61ytx48rKLQri4
8NyJ28D5Apw7JBSWRmGQqkcHKo/3bWL1+ZwXcCIaXXDeaK43HIil9sMz1cZzAHaSPEmV+5TfizaC
yLeA5TMz9W2tNUSVInHFd9/MI0vA8KR3szCmWyRr3YR0NRyfwcdHYYOW8ukHnDn7RDNkBePmPQEM
kTDh629SzyWJpwAJ+CPZcWisxJTeP0ncIdk1No9ktD/c3vC1TjEO/n+oHGcsXwzsS7BRu7H4x5uj
MW3+7Pf6OxjpfyicB7mJKiz9dX0AiggGJvujC8B5HrRlxTqr1NTGtLz24XXR/kf0R+bLP6jwgilE
JYjJSRr49nsssU8WfbMEZLlRxvjf8kIOGUndEdygxHxNQ0rly9IjAuDlOmHzQ1Pt3Uq7CL3nlJ+c
gmM+4+3UoXxwy9P+aiO50VNKKo17W6FgodT53Zpwx3hxDv5jr7bYvsl/012PzY02YJ7iVOVd/nf2
tyBAJYDxPltePPQ/J5Q8++tu/fWIW+8i1xAx+Y3SzkVbGcmKrYftBHbKbJG3YTPAyGGElZytj3Jf
tYVIlehdBp8Joj2Cqcd4gLeS2EvaMi5xGYWun9UBzO5uvaFAdbpN2wYfYlCQI/NplN3plCdbn0HZ
dX57O21ZMPEBAqfQeXdc/67KmSYZiGi1mQmnp2F5QRGMJBG6jfIJq5OaqwP9JXkU86hxkUZhyM5x
SNaIF9jL9pEGGe3LWZAjeGuUM6QGArgniYyydY62V2NVN0x2fgAZmgBQ8fXgZXd2JvtGoHzFPZfX
gU8qgt0bhrZKqMDdwqrTvxsRb/FL+b/oIU6z9MKiaQXgRNPsY7gDktBmieF2pL/E/2PABSU0YKCm
p+8DOB6EDMi2TN9j/ZXMSuKIEeIs9zzTNVL+SiaSh8Thesvvo/qXzFqAUAGavXb9dBy4mxN8HJ2M
wfogMYRvqN+jGvLojo5PurGS8uXby0FefWj2vXXvi1c2XF4h00EDdgsmVWJCCrs01iZF1AQCE3nb
eB7tq7xLIp+odNoYaxfXDvjvfzdA7H2jem34a6it74Zs89Qhjj2lgqmnC9SoS+zvJr6CKtvm3o+/
DBGi0jWA4Sru6kzsjHJycTpzsErqNY68HN+v4xlFOklpCFOYyWiZTZac8dxFLjPCBaCRRqrBoX9W
FaeCra8YB7GYXL5ULEZkfESDwnE8TJIXG8ppf1fVcXPmckgVDgwCFjZKeVYLeL3gym1SpFLiZlJh
Giai9FW9URQEe5fkCfAjVaiZbdLHmcOyN4hN0QEkPjGdNx1sx8BqUUD6HGyXCInSaG8HFaxs7D+6
3CXg0M8w9k0o3QUwoeq9dW2D0zkfrrzXSq+iBnWIawGNiHSEtTmoIWzpzT+W1ydvk8yaPsnslSeL
2U6vOjdK7YsQygfKiRYvG+osnS/C6GdzBgbrDezM4or3zSeC+Yc4UH5dDII4cNv+4jvwVa3EDUja
/nTUA0aYIcFw2eq6iGkmbMsdn+dxvD12yeKMX00w5ZdTOFS16THIy5WI7IHnqzENKnir9BbRf3pD
32LdMCaKyqVrCNrQshQr0gdXbUU4Jhdc9xtpO8ogoIoT6i9MBMVFrNAdbQAETeWY5jPCwZFiSSNn
8nJmtDlsWzugD+pGwLqVeNpmQLQV1UqErLwnZuRLYooNDUC3dWPdHuwJqYcdoQFAojlPcsQKUQZW
GbiFskchpPsS13l3hhCeZ3Ift1w4AYtRPziNwTL1gOJfq//iDJu40tIDOyCIFhceVVBphl5DfK1E
LEshrdWjN96I4Mb7sFWTDttkuoJOLwbsTIT8FHIQxQAPSkBFra/w4kIY8XysGZE/nb/uRpNYyZ88
MVezxtDSMTMGYnsQ4LJLtWkhrYyRsvV/dIxquLUqxJ0Yqe1gtiy7kLEjbMKPgfyMC4fe2EjnQ6GM
7Bw3MPd7asYygz/3Sl9C9uAD92KelEXes9CD5q52M2JW+FqgzlfxocftBNXXliZdIZ/2TNB8GSUh
B5dBuTySv6De1FV+/2/0DaU3M86fuAbzD7JQuovqZDvq2ypjnzQnq2TXF/LK/+Gg8a6F83UKKRWX
sgxm9XLOcWFD0qL95SK2LEVjy2TgJJnDhUeCgIov4FR504qd004xq0SXp2lStk75BlBfRZ5cBLcy
SJ56ZZb0+oRpbM+lZ+qLJ0x2DPDVFnnrnHcoFMNTkRHIcqVvJI7BwM4NY1I2DbNnwEY9NAKVufji
/b3o2ijRypY2G0XNKjqBdLRLnYrNYumUQa0teHLn2VZqG1gm7x1JDEoMw3EdLsSUiMHR7oPhh95f
BQkZL1h0IMvmX7KjItAN/wastOVdZABsm1MbfsCj+c8jZPZcSRFZCyHexTjC3fx12p+/w7Nb4XQs
KN5SiuAySrUPUA0dsH4hstsZwOE9xwuc0ufxTTVu9rdPEHy/LGHW3yKVGHpiVwz/ZVjrfaYCLgA1
S7txJWjMKrjPNAIPgbKuh9HpVJnfTGl0ExMDwAuZpPXxqpb7Id4RTtBrSIGws+bO6GmlX6SflEKH
ATtKBcdVCRAbpMT4yGNxggK/eC3Q+Y958A/XoMIKfZckvW+AtWryXu5VC1ConXQMWS83Z5uv2ia5
kzkaefzTRntQsHH/2rpKWoBR3QEJWvyehxBVwmh4X2H/VVbm3DksaHi3+k4gUGGp5SFN4TwyuQzL
0tx5/UUGIjDns4X3uODXTS4sBMVC4WcPYbLoG3+wmhyvz6iNU9mO8C7Si4gLxRbj1WG4m3fKcTGg
gvxHMN1bNSj+6mc0FXSXNweh4nBy9TbWCAWVE5W8NMOVfxVOWriL+wYc7u6dtk6TWE9HOSlRzdYQ
XMVjXk1w2jRn0yHXQHNKZz9O3/dQjjpd7r4Uag0l9B0Uj/KK9h+hMn1Udc3FdbWZxdiEisGxZmwL
V9hpJhqIsSYS85kdzp1aWUjh17Qf3Kpz+N5V/C3n24nF2EVG0AII/MxMcoJ0NtntUa+a2G3CzdAK
Hl4Gsvhqt8LLz0OARDugexTgEwstHss4QvN98NI9MASCievERl+xgjEWO+288ofG2j9A4V/G+Zwr
5Ewa2eLLtUlkmCIX9NR7PsOFUlTAtqdHGWIxev+289GZZ6sn3iCZ3g3VRyTfaQebrt9MXvCTgva7
o2xOnPvJ0SdkPY7OpipebK9DBfAyQYXHC5v5Bjb+tMPC5UlN86z/Vaq1L3fbyr+ZiE2xhK0MhlG8
2m2g8ZBFQsbokrksyZfcBnuluPxkZ9i5MiUpnSFZPvC2lg3gc2GAJRVWxLS8c5FDtm4MPOpqlWBa
TNZ2YUOn4N3g3Zvv6xDuEZ6Qqj963jAOY/JzQLVl23TAWlYoXS7HFNFWvI2/qQTC/WbGe2HN4Nq7
VzdrDjhP67ugi6REByFx2KRsaTLEmVAq2ABV2qkNRKvMTqFxw7JcGeUmAovdPbjrjGjJ9peubiFt
YaL2RF2CGdgpvelB4VYM7F7rTdsW7HzCG4bQmMxaaBh2BOQcD+2JISo1PrSgGU+tvmVqRq12MuHP
at8kb2tne8xaV27JUruHKeNhPOrS4cXrgwxh3XN/qTzsOIZUUEGfU1Q/mDlKAVzxBD0H1fHNkrRm
UXdlRCHf+JnX4lFes6PAS12sDb7Lvwc5XV95/12L6tRQb2Vy6jl80Zg2lgEexyTNedhM0Eymhy8O
40J4uoc3lt4WGbtQDTbutFrleg4+YWWx6jwsfst1cbRcv8knwb4CQQ8q0xghC1brQ3xoNoB8T7fY
cMpljSkK/Yw0UB99FlXrOd7LeRM4k72WiF++fq4adZrfkYzmdvZDmVt+a8FK7rO9otwHltmraUK/
T2D5joOd/D+xlpmA0jmv2z/FtFuzjqIe+0jlUPWUJY6ibhpJOYSkoyVXDFQHFnJw5+X1J9fAFGUx
RFCarCacDEnWt9BMkwVfsmAXGnS+5AWAEDbYGNnTGbbaLI9TOXMLvYjcP9f4RQBieig/CQkL/wf+
gCniwOHytZa/huVGHMBQmKOPwSkg7pe3Xo7L9NYmYxpAqTr9XV5TqAW9+lHGefsjIDKaCsgtIyAp
VWSIi+irUqgAncORhr3UFbLLy1QUci6rM+uvM5/EpY3P/5DgqUu9KqdBAZCSaywYjk5UvSMbdAv2
kGh77eFAJQ+qkKVzjqCCzi3sXjd+WVqMfu3Pi1ROK/+SvuWuIapqvcxXidLLi/G7rihEVXEoWeUN
609D6vXgl01jGKKj2p2pv3q0RmVaI0xC+d6O8p5aO/lzwR403dNrc7vsYta8ycW/ldG/A4Hvo0Z1
ttPRipKC9Ze38gSb0bxQJIFeVkw8y0HLa0cgezsPxzT0quFVIxq39RWFmwkvawScS0EfbyUnWeTj
KIkJmRJl+ZzMu7qFQ3imrIaCXGtPQxgBG/ZgBPKPSIylyXiCoN31WeD4GohfooW0B14G9etcodkg
nRp8OzfjufXQfRwJzySI967O4G1CnB8dnFGqfJNI/lsQCsS22qdHzMZSLtZYrvm/QNRCYWgT5+8w
v5Hvs/Zeu/oZrQu8ev4Y2ao4QE85mfir6VdhRwAtR+/0XFv906oLXz2cJrxbXXSkFPX2zGMQ19Vp
8BdzW/E0L05V5yDcrwJL1PXwPEggN7DsWhXbFIOam5m/NkMhiDha3F5PkEklyy37wuOhwdugG3he
YER77PEH7rPx9DQ3Eo/GYwVARnes7NmxY7xKuPECBxjIaWzOQG6YEAd4doHCj4/g0xskAnL/+tfC
kppiAgHqDRlMJCeGABIpNnr1IE9oTFdde0bBoHnPuC7FGmPwQSUV2gu9Ed0rzZI0e2xDN/nwerhN
18FDynigrNfVCyPT13cvNSB+EzT8BxUsyZfkBaL/dAKI4E4YsHZIp3FYesDnlUazWVXGMr7eNlta
+qfUUPyORU9YlHorIvn9Mh++Gf06ObDDoiUJcpMWvhSVyt5so1Q1urMvlhTEttLo+kkZQidhShNi
4feno9wq6abDcEc3UQ06s3+xXYs3DpnjHT6uquL27TDR9ZhzMLpDl25pj73fuMkeHoRoh+xE0eWx
yGSnKb2ycAH9VbrkATtWuSFre3vJ7bWkUiA+5zDarfMUNE036/jdP17/xlAIEbljdknWZz9RTzbE
uz8fiT5wMDWul5HiMBN1hWeuTtyljv4hjx8cG72XZJMtc5nuttFCPffN9ISChvqfenLP0274kNHr
HE03H8PM/VgqCk0PF0DJjLPwimMzUcQDVbQVAZz2Yh/saz+jIBp3G0DxK3zWozfmafiznRKgRdq9
FdNBKFxkzQSmgT2J13u/eQJ0aQp/cvPFaW+Xuk2Pst2UDY3LiOpeFNR5zA7KeseWCXbOSZTdsGNH
AhObKVl2xleTR41PqEdNNFujuKzBFLkaUUcSgbbIn4iNyDkY1I5scH7MYafHHztYRRmDW7KFVqEr
oRQG41bNPO5RY/8t15BgleKWqAAEo3RZY/85cgrfcL3OMIQSaEGOaVHKpDnj/Y6RrAUvDOJFPI97
cW88gQCaWuY9RQXdoxBDJazuppSEem/51JQ2hR/bqIvP3qNTGw1QCfOHJ+TmgEQc1037Ksuc33QR
NRpLwIZs9PnfcOQ1GKOu0E5tifl8crJJHU2BdMfiB0zLvwsJuwGyOCtHwkz8ia5v5+UblZQsccW3
W9kTmzvP8GX0ObHP9SvmHicxyYbcnZ/+QjjV55itnBw/k4FGUTCJ/cXDhl3A2xBUxPSf0kh0pDih
GolKUuBGE2eZZWSkW2sh4EzoJbMOglUE/L7sBCGT24N+CARjF7tTRzMS2ymm6lWazky0a6ShV8jp
k5+V1nSdaKw1az02+OjWQrIohYVaEmlHvET+iR8NOyzcRLrsYSjLq1vyXUqH6rjXTS7VejmnJTM2
U7rRA7YhaSzBt1wDIszmzpooIeKC4JPSJCQzSgED6KSgzeATJYoFZrgK7qTheUh+kAvxDda/QHrz
AyyItkdUjoTx+jWkEUVZiSrVHoUdZBlmSrJT0tBBQB1nZhbNYobxHAUztPE6RfRNsmeqjPwTq7X2
2Ssap+0jZpgP1SzFLmRDLHqMSxsv9xlA9CutlAVj5E9bpTeRQzIFkJrpcH88rB45E+rPYXWy9Ki3
UPxE69UesIVnsyGRGLGXGHfKhS3YFHT9KyaVe/Xg7VlMTz8sE40g6pIu8746RsjoK1BLJmKJK0UG
Uc5VDLFS41NZ5NYmgs9m5DkJdgWSNRfI3lu0B4/ux8terOwBf81l7WZRlT7oFIaB/vguXPQRmV7R
N7DwKjMZESkx456hBNOhZgtmjFmTMC/9KhfFdx3RuHWsRHQH3bKLM8zZcMnCBd3aqOivEFQYjqyz
ip/EDv+xlvHctJP9kOktNY5coNn99kI8NEBFvHNEVljB/hP34RJaHxXhyu0kSOBgcX86pnh8I5ZG
tJMYqltL1QPqBig1PCn/toRKQ434rTr6UtGQR1SG2Zf8gbgksV5lj2bkrHVHqC9XGCgQpmcDOePu
9Ei53xqSmG+2lRck+bHIBDD5RErqAuNp0iPV9u93Fr+ajZvayjibncodffUVVhwu0U/ASg3Gv0El
gCwHqyyWJrIJQyw6U7lSw2dVguR7RUplUCNkWBzmGPVHoknq+euCLs3HkliPTw1PVYh5hwotBnZS
EQA1jC17g0lGj7Wd2ky5pM6xEz41tjSEgGPb2yrV70Z28oZpq4iHyul3XUNjAmvL2Y1O0+Z3i7MA
4d1iMVWx0+usGcuAj3eqV0H33tQuppTgfyJzcudlIzlZa1uj+rEcBxalTnKvkHeQzFVP/NGokfI4
7PT7vwen7UqQj7tbQ/92P+68XhBEO4r4t+8BT17Uwl/P3EBUlNPY2qRK9NpeUAKAfKLbHTtrvflL
w75zALMVTQc3RgCSSLr99DtYfBbfq3UQwIlzlgAiM0XF0AcjiU/rVs06atJE/LTeu/RO3XnMYZFc
fFipGofZQFujspwinca0AK9WCu1t3O8ZdPXmBT0wc1RGVHeu+iyv09dgeXOygph7KONusZCsb7e9
zmXaeBRy30VUfvYrvd/2wIe9PWo7tTwnYr+doDXaH5Tsi/31jq9VsA5yZRulZXbNcGyddYWZ7PnF
+LX+5XvJ190Hq+SD/x0/1/AYoY2CEjVu9FjWnV+JDO/wFCHHtyw3Muw41nO5BhVemTnXUJ+KzkVM
68vzgbYdacLgg+vpb0rKqV9NeHHxYAIsyUp/wSnWlnwAMkRSoFkebykUwFJiD9nliXwhx45g8sCR
ayH2RepGQOdXWPNPwnK0moyoUw4z48QRZBXZHSPsPr8rieowl7mS5XFFKiZwWooLVTI8QSdvZ9ub
8F9fZEE+wV6DtI+xi9HOcGdaRKeWLQCskWEzVmCXqn4+6Eydi8S76J76TA+yUadwSLZ1B/wmqj+f
9JdQ78T6RFIDWVl0WxmhG5X5yyf/jWzZsTK2IvUo3zI+IF+NxFk4FABAtWaFvLfnHg4joi3ndVrH
C7ZdxZ5yt0OpzDtduIGkksJ4DwWDd+DMZYANufHlzhE1Ftk2D27bH042kWiWRF4TxfemonS6n++V
vBzvVVOlrUjRiQ3oR633TCBlX896WMs5Sls4pQaBIWY/JJdlfHFk29HYOMIDEJr6HDj6fNo8l3zF
6jz9f0VwatxK9Iw2DEWBKOX4reefVijGAlzfCo7ptubjhMPJO1H75ll/rYcgfc0xVcZVqALOPP4/
JOTwBLNW07CLXFRITZMwCDQOlc3DbR50tmqNnJYuMEyUv0bSaCQS2vNsUNaLjlaj5Jqta/JNQ2+5
kI6FBbOgb04J6YpdVTubrknuzMpFSOnlepKIImV1BBU/PU9JpGNzlKRAfD16K1hwAceche2Y/A9R
ePWOqJS/sHz8VXZqqJXsu1KeQ0yX8r9+qYuTPjR8nwcBzYgnebP73gE29r8Llw9HZnpKCsnro38B
1tT14LMIlxywxXW7YfL4VANWTYkO0tJssT4NWlsMTYCXBEf8CI0/qSGhjp/qWJqLO98hbnj6/q8w
2guRBzhBl0CiCoVTh17zmZ+amegx9fJjd4f5zWvBnfzfDFEEL9NnkGEYLZ4k6jJcA+HDMWn7/dJh
eil84oVNJ1WzhlMtEujC8o/2yU/TAfrlkrkotY0aRcOJmXYgYtE8qJj1BSAUKwXTVzHc2sVqMeUe
47r3WEN3HTTqluo6kA2Tcbn1gEApjwVmAVAftnlAI6AgkolRK31g2bOLmpNLE4YUezhmBksajhWf
dcEZI9AclcYPiqlAv2+XAHPuggzjfXLzFseTv1t0rM1qJTP4lbtC37Mu1UAPBpiP11AKgI2di5n0
8GRK9zfcpIi7Qtv3tVLgew/YMKdSkGBItnii3+3S+fCe/mE0VuBA9UOMd4KCUDl44l6YDulai4RG
frirBGGgE8nG29i+nBUoybor7Yu7Y/z1uOH4B3I5y+wfVvKXjphM0yww8klQMn72fedZ55nMj7zk
9xUnajCm0kBSPchmsaUL+MYKN6jEPjFuRd18jArLhFb1HDjhLmVtiPw4A67ZnKNTUzSgXK35yLk3
mben+fxlKTagf377//9NN/PP7IjQEF7JT5v1uu2R3iL0sRHOr/r8L+1P0q5BTW0U88On5MlugjUo
Yztr2/BvjVFfaWEzRti5sUd2p/Iza7tl+m8D78tzcUYj/pmSB0jGUbmJY6loQyykxawYGKMan/XY
cpRD46iXHO9Kw8Hc5R4agWjDU+CfND/6OKz8IYqYutJz0oxWbO7Q2GvjBiG5GY5+fpch2jr9SpA2
SfDhBftWHC1e2J1f2gvF5weey1A8i4mtY7ykHJ0x8DGPOMZdAb7qpvAwTP2Zk1yPruQoI/onqNyn
TnjaWsczSI142azfEdV1kqZW2tD0KTdu9/RwOGHsKYDirF63GY8CygtseDwcB3xsPEN3hAYbdQvk
i0LHHuwsQxCG/NOBJCG8QtPR6rNsptHrUXjvlTfSr0wr4/GeCaE7+1zvyEJybt2jBrDKBH+5nR6I
Qc7YuqDJwRy4tLdHa9zqiMUTSqgcVtDMsGxnu3Btx9CI4QDAEH0u/6oUUrBtnfPSIGQLHTVGfHQo
ZzXWP30zX3LYuqw6IcTlgsVS//iYq1e2KNGnToPjmchnPxJbTSHBHAgMvSBgnDyKbZzgzDOBuwfr
PIsIJo2s0Apb6LhqnbTd2YVN6cMJUlaJP7QolRzHwWDexAwz0JAY2tai5BZCECUengIB+trva2Qg
qlCEJD3PdVbIFniyxYpWIGkbrcCwbDILCAtB6PTGZYaBXBcbIDBRXdUnvINy1g/HkSdUOv5eGtKX
0Vmx0ZKPp+8szoqt3zbkU58G9Oaf2CyLC2z7Fg9xP5LoGWM0zfFEho28Vk4jJBbJpqNoalhKpCWf
qQlYLiz9QS+6ZEbm3NmPDOuDkHy4Ma/NtRUA/oY3m9/LwEyZSTn7l59PxRrXe1+Vrz6dNsXPYtqQ
eSESdd4AVBZiw1Lhbj1D66Mx3PFIPpqba3+Brkp2qr0KaNyZv/kwhDCE5v0giuPn8NyHKt5i5AaJ
0GdZSRXln2lnIQBrqHsm/DqwN9PlD0eo8JhBZgJ0SgGI035KtJa/1GWz2oD/MvOcIgE1nIMJnrb3
nxscqEwoLqwSI9Y4jKn44cNPmeONj/8npGoTOWLtD1jVqvZfkMWb/pfiSqGT83/JtNcY+dloTYj1
2aLXnWdFCDEPrUsyZh7z37kmDmoYwTYpGCimLaDhxHAIDXS1UVSp4ac+K9a00fKLhum/THDDQ7WY
6d5oFwg5vTrb0A9mjuSsZlWXmeZXI1hJS8gyvyedweSs6fqDJNNFi/co61pMfl++6lX9mlogQQ6d
2kyBaKGGOS/mP8Ma6CFv6wx6GNyYgrRUFjW+72kcy9K97PK9USzh9AVP66R5TIueS3yMr1Mm+wrw
w7b2a/xsmBrfxRob2ItdmeNvn6Ssx2O/NTYVt2j2l03M51mu4+8H2ynOomPymXul8RJPCydtn9xz
6kIcd9MoWYrsgwMLcpW3DOV5NahuIgKxtjIykpwUaOHM9ZKqZHDqNNIV/lUOSu3PD+0Jhn+xhKTP
2eqwvJUmYpa/uAuLWp5Me13wSAjatzsLU6kpv9wji5SM8w1VM47fLAutom8Lg8fSqGP/sWZRyr30
1uRSR2lHTe94/TXvnborVMYj2vK1jH6gL6DXxAX4jB0w3m7+A2c60UQhPweGyx8TOBLKAPJjdKjE
wU2WgfSQp0Xa/bgLMrdVU9PBfEGl9AhHW2wS9jfsQP9gd62wA+A/oRmL1dViH9PLwc6XzuxGfFNp
vTAjxSBwFSfqBz1dJpcwstw0yPujb0MlJrXQ7SFDVVGMCv9yudvWLUVnfAb06uHaTo0xhZzelCC8
TQeY2d7aCF0Jb3HI/qIdgydTf66cjQUjPb92rtc2cwl+uhJLPYv0lBVKxipeJSm+PppT8YmM1f7d
BFQBAMV3EHwfEBW2Poxz/Lo9Oq2LZDEqoOhrRhriHiN48gUq7xVkwvkTSVqLwauabxP6XiTTfiXu
EJ47rtwMyJcaiM9pQUXn9+lvHBK4u7YmQKuWlAasfojl2JUn4SzZ1hAJrcE6yFcopjouNGOr/fHd
LTK9x75IRmOdXcsvSrUQ2Puze7dForSIE4avFhujuaMS3n5qeaxae0mS2P+DtEt5pHfY1Xc/cMSc
TTRCbwYOCMHk4ShHWUwgAt8ztJp9vOUAvhDW+SQVtyy+430tbxzBf/wqVauZ6YZxdpeiPibh3kKW
pbUoKGKGQwt3H4QzKXm95VxZ0NJHP6ltFVTZWTWtGjgCWrk5mk5iOEZnjj+aJk0ckyzkgniUxlBV
sSGK5iXoPjsSh5ambtWIZDgCGojpGLLBuJEJ4Tc2XfVpZBYMTYULWFwXCNLTqIBSmHr0GPKk4xKj
x+fChqUCPCKQ/GO6nIGCOwkS8XGZM2lluQ3J9lUvxrxp0xJkxL/cN/zQWDnef3kYHCPQlJTo7vb8
S9A0lQMHNVVUjDLifog2jDcROyylldGGe6e5RwDygdaCUZerPPgwfPlbnv1m7VZaM2Yt7F38XEWI
R6eZ/iYMsYEF9DQklBQEw19Qd+ffzMx7vIBvqhkz12EqbRBvLt8FveXSlErpKPQanYrNR8iYfkQR
YYCjBMYgEbjZv7cWzFZWWInGZMccpdgVgYOLngObR+D5pcC0EFwSwSV3vwZGceEvspXIk+BQAEXu
rdIajrKinHwUiRTUoUZX99qnpm4Sfa1lpRNIAoBzlGh11bdIViDwlMHRQ+6EbxcgTTMcE1o1tiT+
6x1jAl4z8HMMby1/0vsH3ohVWm044lkZ6e0jeP99z1oJ32EgQ7uAMua0+5dwir3KkCEggPAH+U2E
JMJ1Nf6RnbmK9CZM6Vtg3quRx8j6kx7kL2YgAW2vakon/3LikmH/paF4/1n2JcFUL/XdQAa4EXUE
Mthno0c9B9oMPGCblRHb0Yuz04weqRRZFAVJdPwv+nkpDSuTolxov0jrYb6AXW335eh8anzN1UYS
3nDQ84G5/MutxUq+lXMEsPNiN5dXMclEFJFJzn1b1q6XkgBGAR6FRPm84uuWjIDKGGdW61aUQoHH
PBo0nNU6VKBxO1Uos7blP8+qoppV+ei+NL31oNplLvMPPgd2r81cA5KTkA+1zI/rAkUjwUWoUkPc
Sgz8Ld9++0W+QiWq4u/RcMoEfeLaCGwi3tyBevrO+QYy+XhX03foW39TGLXUixrodwosoJ8KIpUk
ux2ekfVOuf2ETIoK9GxtBdBpbe6ufWOy9jdEoQZ5msrAmsuOWP44dap8y72ud5HS06Q6poLqK45F
KrMe59Vl6YCyq90mlqFXPOadKWFIs/rd6Eckqflh4vY3ocstej87ewHBdlz/T9CVydSiu2DkUsDy
ZAT34ROzEe3kN7YgMlWddscnCYmM4Hz9KGHaYKA/UD5f0dl1oQjwWJ+zBes3WV9FJHr0vZs3THXK
mHA6NmdqhREctIhOwF998tlXcVQXMG027yK/BJbWBLuyMQ8Ypx9CqgQenmrRKTdwgTSZThCbgWOO
+rKvDgmHyyCOiSjabHXdust1dJZZw1/iFBdjXgrARRqFVn1+C0xH2o3lf4mwtJql/Wq5zVYs0541
bBBJP450ZtAGKbenvjrcIWONNnzST87NfFB9slfz4OKZ71DpiYWfXhSNHyqs0qoGPhMwaYbwxlH5
/yuGcJCAGlG5GwwecuhE2CWSdtQD5F7ExzFIPO8VVz+ckywK6qtgUTqhmtzdis++qBYu4xNBy4F5
b02Z8w6jdQUNdwc0JMGHXmvGytW9Kcwfjco6kzQExbbOxEkntZgqlGlwRzCkhSFrCQuuaRe5/n4E
nBOsRK3DWbyQD7C0ygCGN/GMt0R2kCOW2a1wvO2omkRXeVQ2eRytDVLgkyJA3X1l3dSSuEFfynHl
j1oAmdmIHgKUii54/CxSrQONK82EZ9JdeGvp0cEQXT7+XA3NnFpkl1xgV6UApTYWdY90J4/2vtEg
hJSZCLsz6ug1K6HcGvlbflfU1i9y5KmCRavAsX1ECNnYsV9eenSiy+ptXV+iXdlYelCPCdxrDQoZ
1X7DFPnNAHZbV+grBsxdFTXxY2C+w2RlwF90pFHD/tBX+RHBstL/tcLVVvVc89jETYjG4fKJGDZR
f4Lk4A9jF4uvsFPS189/gjZbz/Bo8wH3oPoxkqtbFwYRJC9vCfO+at7kSJKsTaVivkGFuCXCujQM
uYHyJ+FkR49s0bCeE0M3dF8qx+r68DAVOlNg7GUVE1b+eIWL80LgBAJmvYO0QH5qNDe5flylMFGf
C2sHjX3Gtnrshhs1A0uOmjMY1WDkRFtgcke4OzZv8KoKxgjXfgefoWPHZtDr0A7wb+Czu1NNYISj
iamqsrsyQzLSSAOPqJlvbqrrI5mNeMLXdElUui63VasFZesqZ4UqhYHfFgw99iRFaIgtBPR9fKUb
NjL/i5geQVFp9uSMxH0m7SnviS94cX0xYwDiOaR5EWKdD5UtFFwo4MyqKqUfgB7Um9pshhe/Oq1i
lV0B6jji6kruuwCpqgS7ElrnwB3D/tEACiGwFD3ujo0U+Hcx8mcobdz8YyLyOJZ0A9ZW4uLYlycP
DcMoKfAT1O/QkNyZU9e+QBZht/NHpgr/9mqS9gIBld00l4HUJi5DKkiP1h9ml7hkY63Lj2G5qDsi
zICUPm+APXQegTyEQgVTrqMdrJEAYPAUaVWAAisrS6ga4HfbcsDTLV1CLzN0yhQ7ORZjK0C31Lhs
tT6cNOKQPR6pdY8oPW6aCAj+iCq6KP7UtYI7lvNRciFMKQaeuYruesBQ1GZConj/Eb/jzf0Hd2+G
6j7Yg/yM3rNd73MVgmtGLmluGhXPcRpXL4MVEdZOe8c61vq27kbN2nP72lYvMk6RqX+5YoHwI8zD
qlFimAiAlKDm0fwTHeQkzzbKM3SJvzBdIv9lJ6Npgqqdg0sAycmySVSG8rqKWj6kjqHS0eOlW6eO
Plxa7sXJ2JvgtVhbNNE1SFWslvizeqD7ZOSIpiD6smeevmDdElfL5qNOufAeMV+BFtU8CQaKnChr
FfW5hdq7ZOe8JOxBy2piOId463fkzqfbeRra1fIMsG1MAlqdVS+kvFy6Lge8aXURXAy/rMIDW1mc
9UFyY5Q/2+ZMGzbl80mrFkOvNtJW4Zp0eZzpUThynJ+DR00NkJKfqyN1OMeW+68ndZJ9+Vl2bYGF
XFcwOxXKD5HfEU9fkdHjpSzYOUmbB944lEsqaG8MAQkaXGl00V3OSRV1nkyykmDV1ogmA61lJEBj
0z1p9Nbwvb9TCSsP+7dmsPNxUUj4zfh1Xtw8C+KByQRG++SAUbubV3sAdzeR4M7EvsG7g+j/yYzm
GmIeNfQdik40XwGy4Eil+2/A8EW4oGkQcibqQDCzvsgRAV73ILpKOhF0oSFnjWYGx/PDHJ6WvgNB
qRv7RNqoT8LWi31I9kXQ2O0NBXOQ2TiyMH4cwtd7fRViXw2ihoTekSmKq7kQ5aclpPeTCNE3Uxac
iSxcpTFOG2Hh/Iv56+NP0IW9Il/Ylgs3rq2l2pu8qwr4a7hmhpLj9khu5Vk7YNNTmS9NSseUTuHW
l554hs/b+owkX8Q6aouWffTa0AoyyEmzAshKCuHJSLKxuxpXKbw///HRtjspBrvNkbFEH+619Dt8
U1g/a1tlGz4tI5FevyFP/7iqRXRJGy89dCJkHToold3T9GBTQ9+Yv7CXUYaOUWwbsp6HAWDTW4nH
9AWRHaxtfc8Hj+f3pNk9tbBHevGw+6q3g0DHUZBqYwR8/BAWgbtjdZNvo/WgQb6huAB3YEnfvSvi
mEvWed3Hf9bRGSS4kJhT9SV3LxQJcSjDyGJVNjmPC83UNiryD056KS+uiapqHLvqGxCk1w8UgITV
Ae8pkBHNTjTU+lChszi5PQiZMPF5DTYQusQr2PRjkM4I2Xu8vdrlpbqqgJQ5AlHipD4bypDFBwiJ
1LiG23uWUu67zEBt7E/48VYHE17TkhTM5XxTjwWaI0FjAcEx2HSXwe7yqJy4T6lkMWT6bAen6nxK
A3eP0yCqnrX88nn8nyJTjy8MniRSA0BOlEs7AhrHMMxY74o3O8w9o5KxtEQa+yPfrGhZzNwpcXHS
COu+ParTqfablMK10gSo/ObNbWjMssxg5cPxGFsn0mjFpeJVLmuUgp9LXDKeASiEixR9HCWdEGx+
XR1+XIEuwOTvwPMHfCQBG3VOe2TsASEjgC9ojA5bTovh/PITb8Z+0SEfzMMZYrd22EiJlR0uB3l7
Ccx+VVwKRN3Hbr9nPmT+gwEmO5z0IT8HomvTq/lHm+GfHgomyKKZUgGZKOgiAHxemSiSA/oMhBay
16r7tOOp/sjxtAIRu+dkLkQSqecChwSJN2AF4RupP+DhfJQuUqvgAnxgdaihfDAOhFkvpOLgxJmP
QxuQ5LwjND1Xhoi6Qg/Q1nLMG2Ffw2mZGi2nugUHlW3+a/7l9U5EQLjBOyy/tVbwOQeMYdYW4YWF
yFpNabi9zINwoIyCecDLqLCe8X6l/E2xq8IYI6eg3dJpc5/wX6VR6T4P3UwH91X5/JVjNGK2vecG
CoKUlUObj/XscBSBqtOuP3OSusQuJ1tDEl9ImW8+S2yF7UWF50wOS4Z5TcSRS6lMGJ3KC1q9A52+
wylzDw6tuPRa9QetyqETAxhQTNVmA7NWLAcciSEdsIhGgAIjnoJ+281+nPhwQNHYGpPu0DIgH7S9
5YJNkyR5T1Hg4k9u29frvvd1LyPfx7J0VG0Qm6bZqOkrLJNjz3D23oop3DzvOcBKI4/+utddADVL
+BHcHiApfbWqdZSYcTsnwGLIJRtgCGAvJcXvkQaoaF4c9boy8j5m6BET/wl3Bcz9fGnWi4X4kbXs
BAgHKOgCFireFjkT6Wu2ZaexnmT+jQrQUquMM94SDQO25V+6y2XJXJj/eCk4DhRAoGJyIVX72nkc
yhHW8dQnGxABCdafCsvlDTy8EoHhgWv0lZnbYgD6ja5LUohRU9VxOirK5uX/g/tDNuBBAcq4KQm3
UrihkD5ddzLT3Dd59XIvQaazSv79atlRedcmuKe7ARDrZsQPZcYyaPOufCvHPfr8DfSZuZL3+LS2
Xga6G5cIp93SZ2lwdn16yYTVWscarBqjfMHiY9hLTdrNtxFSZW2dSe517ljHU9IsANDn7Ak6FoFT
/8Cpi0DPmnraKlP/L2y2IjlxvI0t2EEzm63l9TnmF8CREAw79skviOvWSNFYM09VBxJZSZxPpoXw
T6OWmxf1E6ZGEcvc43puxIzMExtnM50Oyes3M7B7wm+hXmk7oxx4zYJnceDfv03mCeH+c+Di6kdu
zJjFZ6dHm1opfY6NWtFrZUBaqtdFlRFjULQI7AUnjFx85P6bSPoNAwqVjhHeI2FC2Bslb51wd5By
yinIPYktMM3PGzcLQGKFuIXR/xSbbyOLvImw899VfaYPXoNP5MKN5tGbAzMGNd34hUBxv7tFVYqU
QmZrjTMTQOeXMYCMtJC5qeAkIWuj5RaItdPdqvvdToHXAdzjMugjh4J0Pv9sAV0ho00ZRr70t2+W
GK8L9tP/vu4ZGTgn0CHdtAgHuDCYDGT+RWDyzSjjeyVPSsH5waIepfJBoZbzm/Da5a4brPfxBj3d
CLPdHqMvorG0YXeaIfauOSLaccj/5U+H5i+joTzabrMrxJ9U+1xPFPNxqgH7cI5dxjsqt9nXu1ZK
IB8JPies/jQzpR0jc99NiwGktOr+9c2rmwUU2hrsdOMF0HaRBhmfhpXgS3DUKs76BO0HkjSYKHpv
QX2pJO1xhTo9mvMbeW29G27sPlDPkSbIIMuvSFOJchAxyrVUjLaR7FwnDuTT3vpglrRcrcVkK5pK
sANR1e5WZc96UyYNaYMRZr422S0v2bgKLK6Aw+ubwwmRWc6rfeN1ScOZPg0oG77EsadOizCncZZb
8IwNfVS+OCpWOVdF4d7tbBYi5vpk42McvcqNgkK2LanCawveWRAGTNLusBlZiQu4FHeO21V7F+mK
yL/IQw94+aLZZaTuNA+dwDuX4EoE8iOG33n14OzvbWMJjjPQRSMlgRqRZO4zlwnqdBfEKDG46kA7
KG+4Tzz6sZF7DE52HN5Fi7+iOhlzn7owi4dK13IvZqDExMJOipExOXQ/CSrptN/+gu2IgFvv/E1o
AySh7DpGVgMJ0jDCwsh9xOw9bVgKRqL1qREXoiPUxd8Pm/PpPXArUOAZAyOttZ6uXaykmvMQINQI
czeUxXBKJCIWq4cFnlsu41a81vue5ciZW78GkgERgpo3GeKbZoDfO+okeCVLWW+y29/FuleMOvNJ
/vEUd3flQhHqrq7K5JeLAFQ+CZL5rj/IezGy/cGi3RL4AjSFyt+Nk2Ub2Tz+FaoNH4vRaoldzpLG
74V8Sahs8zfq0jB/h/QrXJo9/VMhaOB3Wi63khcEpNwskRIDn//Ih8BtG2oBbYZZPnRudW/CCl5G
4pg+186Etue7UV6q+09NoMAAG6kYvTMnULaPgipfpPpcB6GVuVdRQyK2KWv+qO6v4F5+IGQ/SiAH
fh8NQbaghnaLu/XUtCMfscKfIgcjNcXjp1fg/is5qiyEyMs25RrWon9921d93Xpsv70u2BJY9otA
dVKVaQvr3wPiKvVEWt9ie5FoHUtXjetS/PTjRmXLRFHp9y8UbtbYH+KXddbGOUhwyhUEArCdc5Bi
tH9jCG+7AVasXjsv5BiNsgaUwL6B3nYCjygYu/GnYJ/w9GTZseJlNLiGwLhhhRLH02OEXnzFXrN+
+TGxVEpPFuDIv9OvMgk2PvRWFOCm92DH+egNgzsOswH58h97Ibpz7/D3Qy6h1bzsv72JIG04Ee+A
6gQcbJGLUuU14KaUBkYkyeSCI+kO3mQWkCEbhvGW5ZCtfJouNmjDkKDgwEtK6L83JA8uBvADHqY9
XD4tmrxsE4QKxr08YLWqvmswR6PKeYG0nRsnqMn/k7YVGi8kIiaDHm5cRsudE9iMNDJIZFq30XcO
w75t+Rr4hhbDUo5hnYD1QikqirD1FpGxvOyB3zK3klkhSYXGex0i9NlqfQj9Thc015M9LnsTI36/
2YFjxE+wWPNAhRd0Ez7NxYh2YoYzq1IpYQbYYD9DXMNFij1O4RRQeImba6X7/NgsQwafiNyv1G8E
1UGLYmvUA2EFgqIyCxBJTZR35lhcskeoKyoGbOxptxdyT2R98nuqOLYMj4PRGcebwLbqaoFLY7Bv
pP9aVwYpSY+vp1S7xCZ1q2ta/ta1xyeIDtSB7LosunH4YvWQyCFTAu2yCnC2I9itFRtBVs64vylK
WZn5cNIaAKOg8UjFLH0KYapMwI2YdJMvuewkKKHn8G1bZngUQ1p/hvsNIfRlVF/7pYJiv79vsi+a
XXQk/GIBBLTP9WiC5QGoe4XJY+t8PAkfWsDQhxLOhXr3Akq8LpUMyJdflBhp9buQavb82nebKLQ7
Nd9kmUZK3qpfF6u0juG/olCz1TXsUbOB6dpP25p2HRKgwZZ+30oih7mJdrFSfgYjHdFMeu2mV47l
0H0BWwaW1xDBGztyYVxH7M4LgM7Ws9e3CS+nCx9MC0pI9IwH9Jcz/fT6dY31evkRrIV3cKpyuxZa
HnNYSu7S8O2JQ47X5YH8ejQHtCt9ovTGluR8wGPXrVs0XWszfuxK3fClyK+dUBq57C7HGUQac2Jm
7GgrduKnB+bjDhwMxRDYHKo79Vtw1vAuuXGD/r8oj+DgqaF+uAnIpVccRlFz7iHvzwuqxWsK7INF
mD4t8eGl80Kr3zmBUvsPAcbDksAftx5KPU1WCg7jSADkoNmQYbFHrH9Bn2k9NgO2hSxiG5IaRdIU
DQPh5q/9RJWmfmK49U6o4grdr7ppc97JdM8oGzJ8WnJ6yE0OVHgLHWnnjbRz2W8d+NMKuPvvX3J8
brsYWDK9FO3bsx/R/1OxHGT8F0Idmoy5psEbAfCCqS3kLwobDzvzYP3K0cXvi4xBnBtI/d7WbfKL
WI6VgYjpyzoiJQTIUYDdBk/U+LM47mtyjQi6jqBEHDEy/LiDg9tQUKWrmC/XkDl7QzVO+VvTeNot
+obmsgV1l0WYnUzkk5UtVFz5BcBZEUtggNG9CDVUIhPK6nferGjXF04Zi2ULfmw2ZuJhbLbdyFXf
6Ab7xczWjN3zkWcSANfsyepUX8ulYOQd0xLSNiZKR1Z6bI/CV+kYGyYUr6Wc+zkRnO/HZU9LbJJ+
jzE7Gonr4JWswm+K+7pkJbM1Q7e81wfSzFiYxhiGV2o5Eb8yoh4KpGdCXuCSDWqA23HOmLAlt9dV
kyG4DIaXkaSshx7ae6KqpnGT26l3yAvlsL3+kI8vaSczZokEoP7RLb83qLtfFTZYiAhOp/r9cOQj
hcWNGhHbZvvsnlf8zcUmIAcWOUeo7XorRmAhTPseCgkiNXyWd5THN0ckTlpPgI0ROQARHWv9vXaj
3SnX0Y6Dmrdh/ZKnjemBfQ6SUTI1T1H3DXLt+/SVuP9LQ5zgd6doJjKZEZ+fzMs/APcCpVIul6EO
oFglA5yIM7urEOoS/D5R11rVJUGBdBc3YXt7dft82jAHpaSE6PzlxqtLHQ6BZ6BWNAiv/goANRJg
TdxSfJbLhfog6P53MTtxkAfdPHXEB/CNS7e7AG/E2GgB2W36xHBqilNm3eo8hYx0y9VnJql651MG
Faprx+TLfmdGb6nco7z0Y8/xlu21pmqDteAWFr0ShtSdhVg/5eoqYPFEhQkGL3fJhKbz7SwbaCmI
3LFD5sbebaVh3OdkFgnEc89R0x3XXv/LI73FsS3i8DsXnR901/OT1AEk4qXHxpC0PibjyXthnZ+M
I8+XhwdW78UQELDmDPY2XYtBJ5waOUlMdeAUOuY+Z3MqrGF4OZWa0lDEHfwlNX5DF04szrdfToGg
QxpGnHuJpDiaY/BsmkBWqycVx46QU95I0DaJ3vb0wHu8pH+/YfGnIkAdiJjUqtqag7jRur6JBY6o
ZkaBgC8Yi6TskuP1fBdTZgWVZw0ANuPdg2pfw/94rm6WBSRtHn4Yp/KTAGYTtVRA1REzASxvY0Re
i7l3oswyS8NGNsIdgXjdDrIflOTuHuaUIKv++cRtvFW4Q36gLCEDcHu9Ou7aRuxObQ9zU7qWuzuA
cI76uIPp83Lqcap+pKO8ha41A/1LvyPIyGg2Tk0g/YI0n/ECAMGjt+5b4GR6or2JiMfDEuxBQc1l
E7nuDeZr77r+Magm030OvRjIYBfcHVDhemGbmyM0SB0jSGvQSd4MXY6y2QUNFcOsSDqgvsjgs0ad
rDvumDnRa6QHjXvTx8HKcTLNmkiOdl00SAvE5YdByEFYXn2RAzBBdAnbslQiKb1ADZzYjn9BBzk+
1N59SWRghYpzH3YPK8d+F/30HOU9bE4asCDl/rvQpwiWMWyCeRZicq+yclwueamHfpIRNLrLotpY
oPobgGJkIruZ8zSGK0F7NuLZMKddLK/dEnW4VkLe7g29uy0CKDjVe2ws6So16hCBIBK/ryKeGtiH
8dGy8/6O4jaAfySaHPtdrlYsIYE3HGJh4d08lsJdTw7Mi2Iid7hsEe4JbIrVu7FB51Ie7+++5COh
D4D5p/op+wrALmorMQVd48BxSMHx6D6U9bNCOisun5zjhIAf2rZollmAvttaWOpKjTqlYY7mFhgW
T9brjnJ+TCcvZorbiEpHbkAkTY++QPvORMdOob2vBhHOQALwX3efyJZ/jH7FH5SgXFLC4Oa+7KHV
ga0yhNTyeE+cNRNDMoxRPG/tBElmHbwi+QdQTHXInHiP+m/mEmkeZQP+6FE8p5B0uzMiagmA3OtQ
3jUymjilmnWX+MEkErRjNQuQ9ZiZw5nddV8R8Z3Rgy1tWK68GuWe9JYnc8wg6+sESe8dmHHV1fwq
MBCwHzzemZJ2wMGZcJjdQVdpJyTJzOuN9X/4kYIWeVcLiOHuq2rOe5ufKHbYK5004f0kVXTY1WNc
pwii54MbPz/wpC9w/B0v5rJLt79Fnu0FQvy3oKUpsFNveoUVwXIcqssgO5u8cTxq+UFdFf6glSwX
zIcxZaDuc8LxylHRt/FeAWPWYDa7dgDb1VRNua1EwwKp6B4I2o5ocXCPBTnPxwmV+j9ZUo8ijyE2
hoJYQu0qdd0k+xKoiBBXcf6ubHCeqPaZVlInZpa2drxsnfj3QLT7Xt5+UaRYS1Q1ma+Eki0d1a+m
EZKty7yiAv5jEdPCOKfFy1MVqXVXQ5apgIflkhMtKpa4FOKwS+T886Ifgw/buWqetJL1RD8kw7Vt
ETUo02TwbpoiGSTIDBIXxkvMb63tzi7V9Z+1msAoMa3iJkUTKfdUKMpFvinA8cU6dhgukNXRCUy2
ycK9P7zGWPkC9JD/Dg7a3HhSnMSbqMPm6rHt/OAlXIbYaz345uOgZvYiwFH1W9ckqFLeoeS9A/Al
SBzRBPWDSDdG4OYqfZCxrskt6aIQTfvdJSIIgrtbpFTFGHNMG5V8Mtx8AeHEkwrtsAJSqbkzxYJB
YvIqM7hN7S8QWIFrE7vB9dnFrAhGaZ5VVWJ7sb6B+y3Vfbj5kEiuFRMwzBk3JqqhS1oZMl3Wivyu
khdhZm/GFf7XMHIF49MqJrK6SEctec8v8h3GhKyMpZ5pn1vQ8q4keuvb5DvmSE2RVQSnuocKa0/f
uUCPilS9W8N87knc2ZPJe7pBrF0ZfPZDt02pm8o1IpHinuj2yfEljkDjx+5rpu7w4ouUMgS9sbUL
DFL5IsGzSRZugbbD0vxNqwkxJvP3powOanjZ0cEYkPBomDp3jezwS8x71qKBCUcRukIyy8pIgHTi
Ac4Dxq3DNiT1iT5gARQn/RNrJYE9Ta4A5v/izDrqhkUuE1bN7Dhi3aFyuQNr2z99wNTLzIpuCynT
qSEU6RcL05D7hxg73F+m4vhms77gR4SgqFU6kC1SdJ0730NnH5F2V2ZySDbclDdNOsW1DewsI5BM
9Rut3tl09TwaSycupIjMyaJxI8uWTwDQQiwxTxXM/qSbS1SpguHrFY37pT653GrXB0B5sRwREo//
h4KohWalHd/gSSsSR6vbjtICgpTUFfH60eelQE+0yTnRv6XzPlZtcuI72U1l0whPMQynUvRnED8R
Cle2S0b8ez6iei3n9+ffJDRB4vL5nVEgww9iZdMOjLnHUVZiIwbHSFKGdk4k7i22d8EUHh2XxN6c
38kWUM9zfdcMWH6fxzdFmfdXExHDm09IvrTM/se2zgTGdHALzisCGOzOs8qVwjiexP+gj97A41Ba
zj4mJpTYZ+gucA5YXebrXJs17vZHDUG/So3afgy+5ZHk+HTExJy8UCVdpzs8E4thDDM6wrMKYgzZ
fcPyrWfZO4G3wgRfV0rd2JdY02fnbTzr+LtfXx0jt5IhvUY2e7g15ef/M2rQTAHZ+yneWgui/Xqc
1IOm0MVj3tH1SFbvhkiub+lZohpe77ctuRlyc51nW1pkoA0n1yufCmXNnbH7V3cvDnIoMD6w4svw
QJsJK0TyHcG6Rhq2QwVtB6bW5HMTeTGIfen8pVNvhLJ9Fj0ANHb3n/wYkfWPbr7XK/wCkNL6/CQk
ZXknrXMg8fZyzKZ44oGhKdu6Uax6anwmVTtnU/eAOl8wq8JHYkbrcL8idRh8qAZUNTVTMojAxOMe
aZ7HhxJYYAY1s4cuZES1EUjuMJlajagEupJjpY8rJuO181pvqknEwazH0w0ggYy89dJ0JAMWOtjY
c5XYxphrx25o/BG369pYcGpik+EtY3Ihc/PZBFM+ObkCgZtMU4EGesN1/Nm122cAOwy/nKm34pc7
MTFyXSxBAUr1G70Eeysh7QcK+vfmNe+UI0w2wP3n2ZyNR8qe4y4TLWgFx0ILsHNqOoaC1/zJv/lj
jexUtiifbQSqBbl7PrZ6D9Hti+XCcOvf8EDrr5dBpr3ioDcmkFtPX4flkvVmQDyTLQ/7vEBUplPA
/fL8B8dabgGgRW7ioLAYu+vcv7SWAa/CqmoomhWI3UYoR8qB0v9aDzGmB9yAtXAhhUTk8RDDUa0Q
G5IoJVz3UXa/OJio95JmnxuAVhDKi0MdRB6ipysoimCbwhiLzX8IgbJxZgiPiAfAqwy+6hkMYHjV
X3g1JlZoyOrkNWm3SeW5VAmUC1XfKNvo/QLngkI7aZTG/WciFWQ3ea/SmLdIwDIYSE9Db+jyS1Pi
aR5ko+Bkyu3Upoj8N4ldiLae7MHeuAXH/b/XdtPMbGlxGrp0QiG78BvTFwcBDX0EBwrsJTtPZKzC
EaUiuM82Yf/b8Vm8/0wqT9k0U73IAjVm8yiM0TTKRbInfnebhnv5vcSvmSRke6Ow2YoEpVRMQ7wI
HwMmNLxnCMi9ab2VYUU1AMsADYDPV0FmMDiy5V4lwuMO3xrYgBoQobMtpGEXVtPEo4N0KRTg5pBd
aRWJlHfUNi6bRoJeiE89PxXhm38HXG4/s+e9roMEMFRQJzby1t/HDmSzHqFJzZ840+POZh/Ua4Q0
JPFhi0CvSsvdulVtBmxM7DTss3a3ypM9V5Zj2/XQ7xkUse7A9HFDdBmsFW+hwbEcDLFLkRJqB0/c
dbwDl7lOX5kTAnOZNBBfNk7edez7ax0tGisjFTZSmoZ+zvKhz5HFZWS8zBWCWVBIZwk0hnx757O+
dGTJb0Q0NW8hxgod4MUZmsQJiG0N7y5U3AelgSwR9d0/OfX++jSTMDQ9CZpec/4ayKy4qn/eLhgx
bX3rBlWhFYVxAfPHm/ZjnU2yj4iOIeJjgtozOcxbpzcNpOVM42CcJ/bOKtvPDvCrK9KdRgzNNoON
XKuz67N6Wzr3r8M3SK9VK53uhTBYpf9PEXTW0c4hUalOcF7vzhZaC3i9CazLYnge3JTQpDjZZ7u8
TKK09+/DSxspIn2KbC9XYdGdTu2mtmAQkVgq2ADSNmTQAgRf1JM+qbRzy6k6e58NrmAQlcWpW2F4
NQoPt0e3+GZPBIGfs6SH+P6PetYz2MCPCK9xf2qMsPzNnPxeGEqGfddze8c0wnOLKuaZyu8uL9r9
DuGuDRY5KCx4jsGgmnG9hsXj07gCS/BHlNd8tnqw6E28eQB1gz2zRc6pI6+9rcjzzhtB0m2jULj4
7nR1jc7JfekDvYweeCy/zOE/rhtrohAJAlOdKVDYdJuWpslmxayzillqYvuyUsIz2N7aNTXFUwWB
qXxFkNWzF113XDWXfC1Gq8f/gxy7AtV8v6qXK1boR4FU9iWAh0p1T8D1s+wuu398HudJkuRJ+e4j
padJRAO7rTddUVztYizlh/3kLQ77Bw6lSNjFaHsYT8GqSLOUS4v+pkKFOUdf/JooYbGdPONijbBZ
3k+50tLqns1GHL9e/+8UFV/R8JwqVrZOQ59l0F7Lz6+N6BqHS1/XmqMnF7b8BsO63m2Is3+P5bfE
RTea6xhnHT7zsnnrwBWZPXLyXHHQYNujjcteMoDPyhWkUBJwzS9Xlxi1FGNafNNQRyZbjidZjP2n
ppUgY6r7TgMpHVXWD4StjT3fZLIaRmKOTgZ7XWvBMGZp6Ag/hpQZbw3di7Qa52XfKB26qfoI6tkh
rImxqSPK/E4vsWZEYP5HAT+/RJjXFc8lUiTJqV2nk75Gecj08qNwVnrV9JU9PcTQWkoaGopGSeZa
79z1ar0qorfGC4VhYpwvyjORDj9ipLiyP2hB2xSey0iFBK1VdglfMG7qu59r1I6Bd/rLYqRDX//I
4gxQvR8CSp/RzNZnvVWA33Z6g+nFKuHktm87NyZzGm/YA3aASpTM3iYSte99B27S9FWRLn5Diua7
0uxmEN9vc4kq81aRUagiedGw8yGeShCh2TxyuMqkxdhVoA8qDffOy6vICu5nxnA8EVWzRDuEDsny
T1jLH8KsIRfxmvZ+zkg5eyTEbXRuU/EYNf69QHIjCzC8eO8/zCH4I+Kpk6tet1rHSccu1qjEy9BN
MLW/O4D/BM3oERwhipp7wgrBIzVY8RkllRdhYmJUYNCLV+gpg8He/9fG+OVOBTqh7mLowCwFTTQI
rArP5Zp1KICsWn6EGI84l0H4pFIPdf25voBOuwu9kuO1XDkFqhRwJfNRjvcQ8P7CipS0N99+oloN
m17Dmd1VGFcLIiKGAsBubEzVuMTvUyFaCCBJD1Q/I7eYfI4QbEL72xBCI19An1UynL7q1Fn6qt1M
fXoiTQ4C0FycDv7xqiwU1jZDH9sTkCHKDS6TRZQkPHiSFxErgU8ZANnimnAhKx4fjWwFfJTEnC6+
sk4bY/My4g8w9pAP4MfYMRDXFRO0sjK0HweFhKWiS+g/vzMxWiyAfNUiio4ORBpARrpYJwVplyNY
BHNt3oIjoEKZPinos3HFSLaGaYhHqPLcfkxGEM3ucaaS/s5iKEZ/l3xR7BaiMT3/5dHM7+2/o4Kn
nIfjYoKFueg81Yw/E9CTgnNqdX1HjV+r6Utp0skbexDKS9fD6Zz+j5kE8/AUrd81CA8kPW+lW+h8
M8smaA65Fhx2HTdtjnyd7C6ND9Bw1aA3FioqA9Wz+HOfLmO9sT2ZvApb6IL+DRAwtsvkEt2UR+ZD
Qb+Df/rF5H06V5biBYpQgrUVvBacnl4tu3rkrjBa7S5gVtVwz9aUCFzUkI8Rqje0luC/JJlAXmRp
68cTh51t+RAqNh2d0M9njxe9D0CbrsLqSL48i5Bcwe3zQscRT7QP0t9BH17iy7aM128GP6bijFZx
cZFis4X4VJMl7Mw/Cuy8WW1OV0uXOnNDb1y/yKB/pU+9/k9EXF2RtyJVvLxaAkC1uSYYt0AWfwib
z6xtKc5xx4FkEErugVn/1gLaVsYcsjsJWeFHoL9YH7q0vjEvYkhyP4PmG4NWdH2UZo/91XmnK4G8
RyMrZHcYY8P5uQdIdZMuT031Usc5DOjJbaHDXyxlcj+eQz/qeNuE0hM8Ip1HL5gKhbVu6RcsJo9U
TvLcdKWI+Z86119EyuDdnhSwWjJ0hjcOL9B0xNbatOhzxVAaCEoJYo9pTTmoaQ8z5VKbMgHn2H93
/Bsrfxthj+jlUlPU55B4rk0A8L5mp+R6GV9OuAqvCp3ksdvmzLQM2KyLJ2OLbnOW1+qsOluPhXs0
EYqneAnpXQkbrRU2EtNrpTAlubkF51kmuLLZCmM6YTLzuZlM+nlhWa01v6wKH5c4z+deot0O+DTt
/XbQLlNTggNuyQHmP+Sc37f4aYlCvaVglTChyo1Ffch04BiDbMc5UP5qTK7l+UWone0mdwiJaF2v
EAUbMLll/YaDpPO/haQfKuI3NXuJ80pjgiGCGHK9KgYnSlWFoM+3trclrUsXITkXrkr2tOKxQJiH
PVi2WxAkj/r9CzKXwpDYi+Si+70dpFF+UpXaaWLyZYYRIPTVvKWZyde/Jz3a0JXbhTn/uC4jpN/w
OK/bkffVSdoMeE8zPvt6gqbmoCH7zMoM/4CZCB8y70RsxNSSKFRDUOjf8r+keTTLfc7zzgC8So3i
axI/IOxHECle2rRPY4Ul05Ca+RlCbvZ7vCQAFn2uXnKynvM0kTJZyO33VfwAuzDUBMoeuPKKH5j3
4nofcELHBM+RZGzFz08ktsMPsFr7KN/GcqjabpAMFSS0lmcpDSpICYvpIHzjj+u+7JSxeIGz/Tlc
duFQRaenDPMr1BIMeZU0LzxrvSJ70+Osg1C0gp1a8fIrjmOqgLVNYpOR4LeOM5Fvl6JVhD+MkA5B
VTzpDFor7qvsfAS3Av50VVx3LcAOq+ReZKO98EgerkDxLw6YzBzb3XGBGE4CkTe8SJnd+UBROVvJ
t3V6uusmmqTznPBM6jNgU3oPihxytNCYgv/uboULS9bgvUSrIRHJqwBatIOtncxGc7BgbRewRkUA
InBXcD1N855AVWyedb6KKhoefXWsQsRnGTO6Ve7z+opIxDTZreiWlLymaJ8o8JVlXoxb2hFgk9rK
yKicGVr4oCQYYhn2RU6YEnCFWeFT1xwcIkfzuEajNXFVGRT+vexy3hPSyDtalai1J1XUolrjw7OR
L+gnIfB+8wWbUw6XeAqXFgs93nyv9KQgP+Z662lk8mx/veP6Rfm8JhmCvKfJHezScl8hyQNCKYwd
DZ/mTX9UKo8QgLp0e8K9BMHD0U2K+XUP06+jGlLvUoRvnEHfXxwc15/B1/dhLFH/KDp50MzKL+4t
WO9u9sjJOSELGa3HMOvzkdw6h2CWRQOR3QEGs5MuT5tcBNUyJ1K0dPT4NkIvbP6pzbaPZ2qlFoHB
4zhgCTxdU5eQQvyzaGa/J04782LQe89Ja4sznX8OXcoEbAHhGxPd8SZmdzI3KGWxB+y9Bf43lPLz
YRizcIUDBWT9d6NgiEB6EwDzSvbrM6b+G07CT3RMwx8YTuSl02Te5b2eH8ivGBkGoly9i12mODN6
f5D7DIypw29qgXXpGsCX9203/xKAZF5TPaS98t8TjIJbmGljWwXOgOr/Z5RRSKaRll56Oto9AQsB
qBMp4SlbQN7pVjKSznqiZcygEGsXRs43Mkgq1vJNDv28nmS3KiNpqJUAGGKskRaQ8QbGz4j6OWPo
jfG2zrSrO6OA2UHSokqb8xMJAqpIKCvjADtXtW69NE1gKxO8d/BJGaZDwb/XH9tVHGXXAYe50s9n
C83D77u+mIcKLO+8ICqWbX6wMLzOfdYJJSaHrtJWSr1depfCW89mU6mceP5HOB0REFvGGYZBqp06
0kiD5q8v8OiuNjqDjn4iuZZiqHQ34ye3+Lqbs44I1rTrKmy1/5kfIfp4j4JRk5hSESu+oHTv8qzA
1l9csOUldV5gw2S5zAkAheh/JYbC4m71BMo8k1E1sIJj7oTK7/EBtNQGOtyCnI30aljM/q8X44FP
4GDf754IgriFc/L3n04xMWVNZKmaM8tJ/CCslQJum97kAso9qGf0WPfRLhPcryjXRQEdSb+lXLQo
R8skiDR6ZJQV/pQ4sTtnVbOi5qfWTJ3BcNnDqYm+tU0/fIPGill0/NLVda5aOc0VthkLwXUhZ+bR
iJcdB3s9obujHRHYAlHbOVYY/jQv841TpPXfYC5c2JuGjRV5zWrwEKZfFG47f/BbglkPr6nVdfhs
evGJqVtPKauoQciAdNo/XgLNTYRYph8Hci4txD+vFIkSN4mJLmpXshjTDnCArER5YBaNlU/vKml+
uRMqMg1JxwytXOHVgJDCFrlY8BpTvpdPiwWLbSJX1ZSK58uECQKcy6J0Qzngnl8jDsXi5ey7hWjq
jW42wQ7f5e6h98oMVGGUg0ZQng0vGGGWCC/SIZrN9169OeU4k9o8Q9vY7BoZ/U+bsEKRv0d8/jaM
hAaxVpzrIPHaDamA0n/uXfH77JNDCYvRtWwWw02/Q+x5yXnLXRvkdO5xGVZfouhcHkG0xLJ6p/Qs
0crDjIysy1ilFQ7JBHEyYJ9vbtdSvQwKTHPFYT2BScHwuxjqtSn+4hEq6DRoC3/YAEkZ1fPABVFk
K6W8FP5x9u7Bn6Psq0PoNnQ7/vnNVQcIgqduLmbuvgEIhIPMtp9Mnx2N9niFZFKOFuEZuDTYFEFX
FuUCAtx4kb7QaykTMzH7T2BoU5wAY9sbIS/8pRWlAWly71QN5yJLdeXXWp0yKZcTRIXSpx95NzMq
ib830mheo3Knx5EoXJY1Bilf3NMdWE3GX+MTB054eav8frfFOiODKyBE7fI9ki56NJWZRKgbthRq
ZUAozn0rfkMvYTpSAFuC+lx7oCCoC+Q6pWTO1pv943k86OqlA/6EQEWswvJPnzT4WJTwyp74gZHq
8d9LsrUJCMo4bEMMCwGC1CA5iPSPdAHIv1ybHu9GUmPFnJgUF07G5FejMBb2cvBOqMgcdR7qxSha
aL6bMvuaAlNlyLY1rRFWAuPJVwUKcdZd8riI/8qhx4UYI2FV+IgmkGc32H/TCEP2PtuATtL48y58
AprepmJCFZNbpB7HwUviu+t0h2XrjXCl6VcPf2rhusAGHPjALfG8t6ErfK4fUS2NVnA4LLBvsiBs
Usz/7qLnxiV2wMdIkxXrWUe50XKtYhVNmrTsdLM7sFUHtR/3+D+e3jRmA+57RgJLp68qPM5VGv36
Q69tc9snmczfKnUDEwH+DCgXfOd4HFvhK/9qI/1FRKsVmNBrI3d+WOa6KhqrYLWjnV18zL/NwLKE
0LYpKBWlzOl2kV/EyPO5RvPvr+FacqY+Y2to5A179WzGqV5LyPmTISNqeCbxhn8iPSYg2B68vgsp
2PF4uJ+pCqVLZM+DeHRTZHB+kFFvTSV5USKnXDIWizmZ/o9ZeKcOSwjS5IJtpIcA6lUeIY3Aknht
pS/PE2Jh3Ly4OCKTs7Ab/t5VuoJsefoH9ypJB+l1M1G9npOYLXLm5IA6+BSglf1nazwxBmYv4mFk
Nr2+EkOTQHOcFjsIXkzcd9COJTLJS3XBZEHMZnkwK/QMV7fLCVAeu4yOi1CHwmZ80VSU8Or7A/Ra
jwdYS7lbRAL+EldOWUDb43hvCDuzlFiMTHTKxiJeAajwUJkkzAJDpfDx+D75JnCrE87i1bnLrUx3
RgowUqrQxSqQ7vDsJrO/SmZgH6fELi7vnzQm0WVXEIA6Ef1jialqcxFl1TIrKshpTz/FCahduFxb
fTpuxMphd9IQ7Ya6chGC0aklFsV8BTjsRMmBEqcXkkoju7BQd70d4svOYABp6K4HyGDB1C4G48zs
uOtLh7IJMWfffhgzJpxVzXE6qcAolAuMUT8UwiKHB6/egNjhKTRf2sjULYxOd+WatmlNNKevkcpD
btn7tqZmlXVvKrrtZDvSB7NjOdekJ5x6IegnsryEWP6x0vNdzu/GU+iWO+EgscdYuftNrnmJXD5O
1J5ibnB0IJ50JIc0FM6/NfiBGTimNPs9wNlbBPC4QhtK3IwQemK6UmKvCZgGgQb7wR9/8u0dQWI8
b3mPH0ZCHM6gaXJ4ujpsp4ZVaOZDAJpgEs5nnPNTpD/RcLQrfRGZMPJkzxHotMZjVSC5eSCfgRoj
6l/Hnw+0N0WHTWuJ7RaRFGBZq1BjyF58ivZ1oexeJ6jDh2J0jjEghdE3pyRepUlklYn7ytTLCacw
7HwAtyyw1bbIvTDSiZ6qjJwsNALFD499v1e5FKEoAnNqq8qgFcFnarcVK4JZlkcoMrNpOyu1+pPP
Vb8VFmie2xH6Ou+99TXoNQidQLcm8MaXKtj8tm2HERIoMT8c0WYo6Q5yC0Mtu/YJis2rX5bX2iLW
Wretrf5bjVpJUvygl0bU16Aw3KzHkPuTMIL0SAovjzyajpeud93foc5uoz6LIpJETED6GM99VfjH
+i7qRRAb25cwMtmq2BtEChyBf/4RkwKnIdsNS8jSemCbvbCGhzlVRYHwCqYOcDr0+FsvyjaolQny
8jMBvkTcEFbolmzndUdy7fJDRQnT4vfsH7HhDoXkms+6bkbZ7FsPZoSA0bL5qtJl9LNPdKIAS3xQ
1ONCab3bAtkp+3FWH7vsMSfXXp4c/3H8C/wC+sne0Jhoosmt8/1O/hq4yhWJMc/CrASXHaQt42f3
toQtv7N+8spKWJ1RwrUUFlRptIb8xRdORy/8MWQPC999bI0XcACCfmdQf/2OMwfYER3huEZthjB8
OgKDmmqzPeh+NRy6ahp/AKmaj3OWpjudbZdrgOjHVsjjSty13U6FIB61Yub0Swxy+dbE3PWQ3zsH
BPUFUiG48lnz18W/3jj/kkkBPUDzB//AxAqieMyscXutyjA3hEMaqqtoMhf4NJUkspKGzHs6ghNx
NzxO6FWi1BMSOTwQlBnyzFq/S+lglyqw883LMoinmmnwekcPzut8+og6BvXF9j2x3G2YwnIsr8cS
QVIA0Suwgdw2+67w/ptCoKFcogIPbiWAbHw3xw/z8QT+uy4zenR6We0lDHc/ScBNsHPLILv11OUr
g8UzOo2Bh+NAnAvBnbTlWVxYtkAPPmDRhd8oTID0tbb34e2Rmxc5oxqp8+SwlGaoK53si3w4UnUh
EeQFbcSUqHuloGx7NQEco6lGNL6phn3oTGHBzCoU1+9ddnGvTvLLLi6JfAk0r4K3Gs43v6yvQkoo
vDNyzmg4jyEjLs0sGMZ4ACgKKkYGdVcC9N/tmdccmiTZBLAMkXbHa6XbjJo3nlKgfpbSYBVAMVBl
g+0EHgCoIjMQWSoVk71UmpYjtORq+bMnQEk5W7owZRGemYSvZHzAXH933AYhQu9PXCFgwYwgTTLj
aCM0Qj5Jl/Lb2Sv8wZlZQkkEgvasCTZu2GW9N3bmbt3hmVpgLlUJ2rjHkCJdKbZjyws4Y/sj+g+D
gGCwUpLOKIBTjDOkw+AXAcGp+Mje16CeqE+oU8VEbgrP3qfTywTr3rnEANnqgC/LLsvG0n5nJNu4
UdeBwG5UEzsGIokk71nBYi0D0BCZ2E7g42Cg6pciVSP1yeesiYeZR8Rw16yWLKoPHFPA2y/pWOzw
t8vqkL0N3rtWPCTvjL2mROLwc/JnLBHGP4XW6sPqE9wnqu9hXFny3szEJa1XNpXY60tmqyRiO2sk
Qcm4zxU3dkcHSekzTWbfBwAJSRqdDtIfjg6JAN7jBFoR6P7cTHJZnvUwTB0m7Iu0VrCEZvYZyIqC
jKhhhzMpp72KzpjJ6dLWTX6cRPc1kW7EmdGt4ssqiGlf3SkpQjfVhckhqOqReVonC8243UsBTTYT
9UqpZKL+ZsbKhNOULHyFuXk/tCDok2zcNF9CHi7l9WNJdLsX0mdkVtnPzt43SrxIN1LrF4OV8aSN
BhGLRlG7Q7bQTUhhMT9GF3/iUazrDgf9jcT9rMKmeP5AZnRpZ4otAq3aHfvuKgvddsADzhX4CnCw
h0MSpilMuNhJXsuK2FLMOuHYl08hefKmEkPIxY6Rr3s8Wp59r0bnGRLo9tyUO3cAG+lqP+aqhtD1
fifPB3G5VUDfRRSg6KteTCbBMbiHPYlsjIY2smLCilShwc7Ae3/Iu8zbclVbgWCjteplf8DCR1TF
t5bldkbsTMwu+6bGtjcXXFc2vtAn3oPv+jge1M2qZapysHOvu9cwjBxil5y3zqvv8YvdkCJe4SZT
u44Vp2EkQPGscykT+ZV3LA84gUyHaGpvNnhkHuNuYEdufK/k58Yq8tOQm+KYsjnff34gezShFooz
o10lmd58CD1Erygz0IQ6A9H/yX4flBJo4Uw1/epJ9v150Rqnh/TErhhQMpmrPytr0Nc5jgYzu7W6
BD4iEOb3ACn/hQ5bKMPLhdmm4rYnbGhmUcpn710WZAvUkXeYrUQbJsyX+nIHMzfwZW/bDb+tjAg8
4bHSP1d1Cag5uHih/E8IZSS9NWYwEQXTlxNW1X1Ao/fdzBQFEoDAjyWTLgdFNXCYR78qKKtSmRLQ
6236xYl32oCC+V0sG15kGbjwx4GMtj1jenQwIj4ZDgLyvWJ/bniTigskepX0fZv3AdDNty8JJEO7
QACTLZsHe6pv6fhdK5DB/GgRGCd/P8LvsLlSaPSEh7vOKtkP4WT8gWaGfYyCoReeEE3uvx8fVNz7
4tlXQ1LgZ77LTJYQo2ETtKa/LqkZtPBsD8wWruHMW7kavgJ0LV63pF4mnfGZMVf0D53+2jlxZfn3
EV659Xc6S7pq7tO6omGxZ19kr/uZTs7/B22hRlXTIPZwm8FNdZCylP32/urMN6df90CSaWXoUDue
E3dMM4YwcWZYE7wbcfrmDLCxLYtCVnJnqoil/x5R1PFm4LDgFcTzujUQH3Sr00ePWZX4k8/QGa+i
NzjRIAdwydOxm7y0PwaLcQOfdOKDZ0eVjxkLmMrmYcSK9my1vI9ZvWb0oPdrmPK4F17Yh7qPdZGH
LNjjzTFvKI2m4Y8aGVoo6zKHKPOfBi6xdU7DBkHJIhwE7HAZ+9Tn+fouc4DLxGa0GriTdPTnHy1Z
lM+bKCeHrnWv4iRnNofdJn/+bJxTCXgPD4xyPLVR2yVfEDMedc0awfWyA5w3iNTaZQHsftcP5d0u
qij3gmLMvFjLRx6oSTFBtLiyb2zhvnjk7IqDvpGw7UmINv/9is6a035C9+w/LdI+pajXYtP4mEyo
zdfJZjf8B2l5kqHz3g52v1slGz9FbkFNFDYrXlGfkflEctFVXNjpg6JAXmo33urGSBf1u1b4/9u3
Mlpb0b8Y20PVNNhamEIwFK4VriaDfyajfeclu33jrTTJvWfFVM6iyuA/vQE7nLhOaUwU3oa51Naq
btfMb5aXFo1fCJP/yruR/fd2n2tusvn54vc8oZgDWREH3G/oU8Pu4jYG495/S7YmJ1m1FUOsFa82
P3x7m9stEkwsBQFMKAzJt9764iH1RHMX+Tt83AOHO4q/YkRl6N5fkt0LCV86kLiyMiNqCohIlD2R
dynAWNJK1l/WIEUl8vLoGCNCOvWWTmhIJGYEWENi1fU3GSAf7RO9T8k9uSLdXSgYZrbtAbzzrkPR
EpLtHhmsFQUHYfAXvNA4fsBw0T0tL1O/A6tEj5KFyFXRgD0o2cs25ekAjnYoUD9/a0fwBMBQhWR+
18mCyvRAiHORlVmapK8pinURO6AOnToySBLeTz17/F0ZnLhAaOFFymO/bb0RTa4fK6cWrdpEALib
91CLzgt3AV+LsrZr8TjL/shQnd9oAESHM0AHcdWCdWXcsZZLAXJebS1W/Lg1N0iHO8Ed65W5rK1Z
6MU1COZuIAduvUG/Hx+sJmY6KOHUU47TrjLy0TRXa/7MIyfUMJ7o34KEtIX1pDQCHXA6yGel4Wb7
xVSHxk19HzzAu0VbjN/vu+WPQOvjcKO5rkZrwiYcjHkXZ1+BrpZP42n/VyWr+v8CxX2QTXC49fwk
sdkegcnF9dJ9Jl44mlOMT6C2pIgUmf9wfZTqJ+VMwj0a1Zw+r+QjlXKHQRxcmf8cyv76mhb3kweB
BsPeDg3QwiIwhggvS5h4EKS2X7Coa8OuL6UgyaGiMJsIpi1xkEBiWmv+hhqxRe15wtJfiE81EJb4
IhrjSNoSN7SuZBSc0FUXY+m3hXmql9p7bAd8lJx3a2vxoImANiihPWpxNpleEKa07QtYchyaZ9uY
xT026tNJVaODSSXwl59B3VmtLnQwW3h5hczjN6yPiYPEsm6a4Z64+XMWans+vgJLpyHGRDlLTae8
ggFoc5NDbcRhV2Db3EXh3qyEGRZwTLjX1jULiF/ytUdkC92j+cWTPAOfTU+p0NwbreRIjpMlttXo
8C2I0G37ZiMOAztCGe8KQdI4YF29i7gDhatW4lRZygFbDCIgNzwMJtPqtc+ifENkyhsLpn8Cc1+h
+LcpdIwi9Ilp8Zo0NPxoU1MLbRNuERfv6E6cpYGEJNMeUpGq4yC0wU06g0oVGCdCII2TqlB1SDLB
w6z7RnSMSfiedbRtHFjChS6e2AnGgRFwMzUPEmuz6ChPC1yCREa7r1vEa3u/Y5QGH+b7ZnXhu7FQ
OkHuA40SbRnvLA1h8SjqNHsoVzZC2QPzWBt/wQ6fktT2ZMvu+2ksyOyOvM0Mk7F1b8Asuo03EtcH
RFTgbxZESq38v/fNCW+/eygF/q6yOQMKuAlcg45KG10O5mJ8ihA2wI6P/8cgmuuNGehzjSLoJVEO
b4l9OUXRUPDNrTG4GeS7twp1UKOBOSzfd1iyz0x2MfLmrbtwGqbN3QOktZXgAcIM5COQ8LvZ3WL1
VRhNSuA5JOxmls1jPPNEWP7UnvX/qSPZZIqQWqnNSJFttgN3+wV+P5PQ5Z4xwc6Ift8BPGD5LytS
nQttvoh4MQQ08oDmCAPpJ8uNHWUx8BR/IsgKLqfA73MjpDlFfj6UNAYLKlQo7IJbem7cvzAL9tE+
Q3n/VzatnyZUjwiGPjke+Nc93uumc1gZhAy2nzYmLVGa/s1AILpC0uYKe90w7Mj/YyegeU31Uwf7
fm84FTonSooNjSJfhD0mJEWk1fe5iUgKhC5E6RGw2l7cbLuWGEIVjoJUmZB3XQ4UADXRA+xk6jrE
kKRhKAZvDTdaxsszUV9McdtmztujDETOA2/LWcSjVvqrq6Jsl697UGr3JSdDlhPl/zga2+UczLyq
+lgGy4vu7oHBubvh9HTdRolBO6op9Naf1saRKx6z4spfHj9nCf/OVguFp/SqLiwV5Aq/OAt3g/xa
v285fp+dnBrNdsdDXLI6qYcDwMnIXVFHs5Xa+aU8sMPR4O6Sv6X/UtGtnh96LU2/foIAiox6yMCZ
cXTXvP5D6hZClADENovi5Knhsk0KrNkOm1Tat3XRiB7hGkdLBYbt33EWgbNk97JmhOUDyGAdalqy
0B3OaNpt6NDRyQaFHgnEyxIH/FKfB0wl4VIrMF69p2qtXLaE0Bo7yV1wNAQOFU6lrv/iFPaD59hJ
10e254TQlGG9ixaCs8ABQ/e+p3gjd8PzDM1WphPRvtkrBPS/tL8/W3uAZVMYKKfQ/hKK94bXbJq9
xlcvoQVySxjto/blLS61BOrqI1glfVwGDzI/AvtS7bXg7nyeAqYyUW8iCCusqNclyH4nq6SESJ0K
pkBWQMqewQBJiBnj5NNvPga1M6E9qIhbkRSKggavH/Orv+sDpb14aWDqZNJsO1oa4SZPSlQDGmk+
H2LagcmYLbDpGEiWSk551dJ0xozKCKCp0TSfL96/9PzZZ2fR5lyQxWRe1jQPhPqBwKci6DjFtF/y
HqeNkepzpzHV+uyII052NXfgg8n5AAclnH8f2Xvpgo5x72IUVogBsA6FU6Otg9vfyOCAwCMJL7QY
JaqM6ZuMHUHe1FNqnumwQigGJStg9/vR+yrTkwNoInGJffS7+EVBeVp5E8SxsFqT250dtCrdBapK
Nr/384U0MQQrJ27e+Se6Sy4ZMwcd6B/8or9wh6DIz6JsqFbqwPqvquc+zK/XG4cEgaDJIgpN9Mrt
12ntuPUvn72micYrT3m341u5kp97+wgLLAyTF6j2MSs9X5Zl1Cmp6+mA0LdXPGfBvI2J+7zNnnBa
aFLhu0tMZUCJlXNUK9q1glZkyEiJC/1bZQEGk6yBLYiJwYjIaUctgGh0IS1pxBl9y60ONRWcNukE
/vfj+LlJ1lcAMVZs9MoDnuqUnuZ3YAAWh+kYWrvmoBzig9bmqmykbMha/vc0cDUw8+7ooO6oWPrY
fFU7oN4zs5XOQBqyYCQt00sEaaVsrPbs7uZgFGsCKlgEhJGZI0JDMHZg/B0YDoizuKxwL/3G1J4F
+jYR63uSb0BBvb2DE3x1sMbjFuqRtnwT+yw54OgO6aEh67Ue1u1sk5KPjG1F2N22c/8bLjOzad5A
sAYVJKsOGgiARdxpt3IvZvxKyrIo1nj+NiXVmsMI0stWE8IA6q6fGsSi2tiQe+Mp0TZLJvt+hOZn
ijHxrJmEzmGJYg+7fKp91JNoZ3xvqGJaIfVKPFExx0qZaUWyo9TOrmMxa/JZs/suDURZXUMczEO7
7NqOO8+UuHSMptO03nAukg5BepdKNP5KeDVEpxoPMaCBI+P6KYiOiJhMET/M3lVylEXUOOdetybm
Javu8k3qQkZVw551CKaI7HBSXl4yjBJ09N/3Ja2/6RU1lGcSthNrMlUsQmqevN/a+7R9i1Z8zWgt
7iZbzbLBriwlnREM/kdjXuILL+0P2/McfurTfKpiGS4aKfzI355hCD1qEtii7il+UOyMvqrKZMGL
HOij/eL2SmAJGgZY7bcqFpeshLGtaMz/LTiL32/ZzBdp5A2gvH7GIOmqrwED/xgBsHzerilbz+ha
qwKwaFEuf5hgkF94NfZrBUKvuI9AKrlzcrGc51zsVbWk7jVXBHg+hSs6PCxL65Oy+1e6Bjd4s+LM
uXx8xGcrmO4GLpkMcUeOcZ7kP9XVpTlwxkTPQrzxsfBcw2JTMEnxTIHHHrfHwp/mOreI2aP5/4l9
LSNbqSydY8pBuBHBmjFdVVjW471tkjVRQJPro9MoGLyJzXDQj+vyNIr5n9M7BV0Zauymr/Q0cr4i
oznXVLa0obPvkE32tsA/eG7AY7A2jGPASzQLlIYQuJilWerztg9R3uk3LW/qym3Tsqx7TeMN/h/w
yAzGCTTApp8HTJU0VSiLA1Kxsnkgt0GmDa9G29UqKK2q17CRVrEU43/vwCDnuU4h8Z5pzMYDulfr
dLxVwwRojWM15iPNqiIqS8dtYZAqIBFuGg3blujH9oIrW0RquaTUGnB4V8NIi29IMXSRHTjZn6YK
9vdbkgkunQ8R+Rxm4LLpRQcn6qhSO2eIE5J1IjILGR6NdWFZyNvoOMw2+Eur62Exy70m4X6WvEat
duDtqMFv1i6wXMYv1DUDj4to7IBB/cAWRwgu7VW67NqqDsshHo/09728JG3ZKrdxNLoKbSMscFJ2
4zN9c8tPH+nbyaN9XIDwaXLUZWN2AzISR3mwRbCCFsZmKeq/nnrXT88My9UtVez6eaG7hkGaK5eL
Pmvr/4QHo6g+3gH5y/ej/dY+ZC5xxK9JFNdctmJUoGW8yW/hkDLRhx2PyY5oEkv2i6IeM283zP0r
0XcTfGkNdwbaMK5OxP7QQmOuG+XdsS2gz3wL5+4xVIo+dwR9w94wbvgtwNaOTRYYGYTQYkeRYNkV
CVrbN+3iD5Dt7sUMwh5lhWo1e9SVohLWT/5EJuuZYwQlGrZptQZ8g7Wbu52fQ586kk4OL6rrYPeu
Yj7z8ERTR5rTHq6mbKdJG/4nJW08+U1PEwKkTLat3J+WUc6xUDj7p7MbT5ZKw+0amVt0RFEmIskx
s3GUrwqQjB02ORUrPR8i/UiIA7K3Nhv9URzczhh58brTjvqNlJn5U8895dR2MB/ewimi1QgXpAkf
Sc2TFXvq75f/IBtwGv/LOxPppQZkIbDSBudYcFKMwxMFonF1wotzj40M+bM40EZXjlnrrD75hTvu
6U6yNvNf6KCFT+L27R5Sodzja8l9Ik3+F3WPEeXz1vCOA1U583kFaoRZjCmUm5EpNU2DEdYMb5lv
UA8YYWTNlBfdm8b/+91Gx6bguJBNwqJ4XqTuJ/MoLSpRQgfplFL5SIx0CbRBG1+EmDRCNsScCL1V
VqELwWTYGB6l7L00bX7nSW5uGgAgaC4Gn9l1KMfh1uyF5hWiXhuslsdqkINEvFGT7pX/+8oCw8qr
dfMZi9RU89DaW1xGXHiRtmKjPATorTFbDks6v2wBgT5unyN5QfZ3hBEqjDU7jmJPQfTlp1LyoNpz
qHXF4RzMKlohueR78lAB5rHuyxUTLMi18A++E1FelATO66k7E0k+sOySI9EeZpwe58Zgxzuu3SXo
ykYDyyX54/Jtp0BJXnBop1B0Bv2DdoHpc60I/VuHN3udqmtbYwitMD1SYf9buGpI/YNm4EJ/uFig
lU5hVEtIbutemKuULcY5Mw6GNBvidsgiUlO/Il3ANiP98wU+TmcMEGIr2L2f0kddYPsfumARPzxS
/YOrT3NW8JLEH7SLF253lDlNNeRGz3ZXzv50k0TyWbgnOxXQH5/yMEfPAAjsUpeMGzjASPLXQYR2
gPUHRYDU97J8L6J3MM6EiAwhhB0h0xeoIVyrvZp0Gqrd0X+sO3akCovcsrRrRDfhiGO3OT5ubSZy
tFFUylqbQH8yHIewlLwg0+E7viTYAX26W+SMRkzoBbk2bgCipJEF/5/b0A6/cliCJKMXKY1j6eTL
AtT76jkJAadc2zhK+MsSH5pEaH0dTu3ZkaMpI+ukqEwmn1beYrFza6y/F2Ueyv9a7a6nSX/kFZCZ
qhlUiXZEIrWR+LX1MiuZddCFfEzsJITcdlz6b9EoJlE0FzXr4hJd+4TRYnKreJQFCbgpK+nWcKTM
rPujXfptVtK983z9Z79ZzQeEWqG/Q91vaa+JS51O1H8xwkzzR8qjQIOEZxUQf+UG/ih7uDg8RUdF
6hbvUDruu5izvIWRc4dipi8WlNOLvPp8E4Lu5b2VqL/zOpjT0WOcs5JPHIbY/UKEaGFDNKfyChZY
4p4AlHoZpaZ/y0y4CCFZd4Xpne/koRu8P8eYJjwcLKwt3sY0w56C14uVSDkOw/QNGSlOpbMrP9P6
V/xj9QjRW2J+O2e3tQJlZlW7MHxe6xp1AQksc0SaTSkY6nEZDmbpJd8AiZ6feKuufZvH1y9a7UZL
80qVNxDenG2zU0J2uG+uVd7vO2lK/Rekw9UdZaZpk+DFYpYtqXgEnMp0OmRLUzi5eH3ioZLzVzIq
uOBgLV2Uw9M3ddjjh9+AZ56qktvbjfjyh9ndJKXXm1i1/pnnuJLIHP411zJW8tFhI8BiMRMIsflV
tpS+5bbGytF3Gh635Z8kmVN79aeycqGMOxh4s9wI7NnWFX5YawOqm6JfDctBOW5etsO7qxihL1Fs
DHKiQrnTr8iGoS0+6nL0wqcG4s2nGfw1MPan2UQ/E5XoGDtPvrPsrfOIiVnhT4YY83hAxzysAiGj
q+rjbsY/KBdXvWt6QFArwIIvjhP5tLmNoBJDO6wfM5bNx4HYDO/Ge5jCfJbynkFLMmDUHV/Jh9jE
zpWUsLlo+OWQgQNAL0hXjQeQzEn/ZIt4kMkub+1Ntrj6R1GgvopXvExj9mIBUvYaAA+JC/tQ/JBn
p70RhpD0x2XLBbQPzMHjIEu3UAsoFLycP3G90CJ0kDjRaMs8wlbRWj6EdMdHJJt77MgJljkmBu52
VXrEEmHKKkvqN5GEq8Xk2u2y19CxrmXc0/M2wioMfriVTJpkECVOFD1C8s+7Lhg7gjfYxouUkBYq
Iw2ShgoTYx26bYFdHxVJtaMSjqkZPnrwchUzyiE/vYYUbCWQGdB0UJ9fRUpjwahVfX1r5Why2HRH
o+SAEHe54LIqK7nU+RwjK74eFVSMlviGAvVrFQSKizqlWn1GKmfKt3PDhf1tIWZLEto0+nVgEQRe
uysmz90o0KqcVz/3IhvWOy+flz+kPeLiHqUjr6Bye6GA5OxJNM7t+6dds5augmdxIshe2y07XxJG
OND1qqswD2ohQ4dFMVt5xr2Kdi8Hul3SVlQYvdUda49clduUolMRT06MQFvzWNp70Awy8GMiLQuR
aIxVDddSV4n6rZSMoZWx7/CyNaok6jHX4C4jzRsJuBOE8afnswBreA6rHGBsa1r4utdM7O72b4x7
ccHC+aM7TXr5ye5lVtMlv4gDald53pJuAuhaFjTWg7lHLRP7OjmOMntNhyWF8Cnw0UHoyd3PmcMF
LSG8v/B0t0c5QpSG9ipYphXHTqcbZEP45S3GsAWjPT5orTSV+fawLPeu/8tV6lunfraTJMdEDvT+
sFpyYD8H/VqzgLzOjzbkGJ9IqkkmI8iZV1HBkK8e0p8Bx1E46NNiR4W8SRnUxXJPZpx3FSZngItY
BRdxPYX7okvu9z50SqbW4/wuRNaq7UUyOwW2Yu2YMIsGWCzwIKkyoapzS9N5TlCwsrBXrzh0qKB7
qYYDwfQhVO3bn/qP8sHLLQ4hyczkPHZKt7Kz5z8zNUi7Je6jZGzgWCmLOYYvT6ZjO6tbhOVaSCv8
Qz8B70hNKFx6M/rkJfsuS/8PMJLXUsNu0iqZ/tZr1OndOsbY53CrajNHHIxFXiLZ0OQfLWFUFqgS
xUJUDtLAcKC6BnRrIhC0QvzhFVZvrAzwvhKiRFw1wdPKQnZe85cW1LWgjfar8NWA+lIgV6L0CWo4
c2oLoxhN4umYSLCZWZogFzWFf7/nIlRpHFwAYkPBHHkLNSL/rV0MOe/+DrPkQWHLi7vrW2OTxxUz
xOYXgODfWRHZSMiNLTuadqLEQ13CBGUIT5li5mpN/rgx6E9r0dPymb4B23lgYzAOoM7Vic9tnycx
2HwVQSzDGz+0UK5qrYIfIkP2HGLv2hUO6salJ0MU+RE/NfGANqqL4XQE4CWzgpSgfieehW1cu8Hy
HOHj/6LYnDSoGBn2pPy0qo7DFIPknmSCNKbM0rvyTA2ZhWlsHPhj4PH0tLn2wWF3yRDG2f3F/h8O
qWYpijZqes0HNX7s9o0VVmLkzsxCy2VevjacXwbK3ipvxSzgOR7mqJtJFYtsvnKocjnVCdH5ByCs
9vmO6DTOoT4l0VyqtrrKsfciwmR7gJEUPQknDaqzXmC0yhqjwsJsqdY3IUQ387cXuuhI4uPunsDj
Coha8Owl/Y2TH2/Lo+N/yrXicU8HcFI4PPwkHz1WriuHFiMBUqaDRDZ5UfipJkBEZTmitOo8F7HY
0o+yU62kfOIXy7+l42fQj/R8oAmUS4C0d2+5e0+m1SU0mjl3jERdp+eIog/mu9DIpYapKcuBmEhx
95R4WLavkYvpVNKPztSXCd3D0H3a50PTk+nkzaQ5qyrcWimtNLy/1iQxmhPp/6NK2M7E44qxQTkC
p9tQfG2s2uamoSqHpNzPxFuURcWHqcmob7SROInyrE1ZD7FRsQ5ZOpyczufz9+qRvV3h0se4fySS
EeG2muuZ0Rbv0SfBmYA6EWewLavrE4FpVYaYvtgXLhr9n2snCBQRhsg5eCWN2XGu1YRN8Lumr+N+
WcMek54iXHz8juD6w1zhszn+ShFsWRbrjUSH9OKC7MTs75UBu6wg4aUOdIpXY1sbSr+bQomUgY4o
2ikyeYrhykZsRO0ho9EqLGs1bBhbMYvp2Sza55wKe5gBiTsOsNxzuxiNRSXl4CSVsLJpdpell9xb
eNgicD4yjjFAo11+qRXiU9TjVy6OKysVmK77nSmkQpf0fflzkbtspLGoT2ExHTVwavvCF2E92ZOJ
OXU+HCVK4OWoTXAWprkqxj9rg/zlpc547f2I1UJG9PaXRIrOHy/TSoIcXGOuSt7UtlYOQZWGqDiO
L96G8gt7N2Kx9lIObj1NvO4kn0FJdP4EZe4AFMP3DhleFVS4ffESiWIryxbGnKx7HTue+pbV0fIV
GmNH4lZ91lxl9WXD/ci21WAmBsfwgSWUB8Ks3JZ2ioi7NCsKlzkBsvt9RqHYzdUpImw5pKUtQvwB
aDvcUr74QNeQVyt0nWidaQoVtIkSQaT3rIA8nGAbU40m5D1zyuyetm2pc/CL8F0OlDBhRwCTucl/
yIiaphMfDAyPE4WmBoJg+JvSkZ5EpOwlq29Qeubo51z0/WPeN/VJci9SbPtXFpwE0lR8FN7M3gmx
g1KEMU4hNOfyrkJ5queib82++HqPpjkjRurbc/p2pLYjU2gH0EgwsSTDx21bUvUNxiG4e7ROfYo0
N37dDZ1riLzIi43NS9C7uq3cz1YSJ+P2eut4NZ9fdI6IiNyctT+LjDQxwfTztCt8R5qQYNHsYqzw
Zv5vZUbSFCUcdULqyGvzVh6hFdYyHKHO66wx6K3uYS+B37NhVN+qHfHffxWyWIXDKaM0NmZG5n8x
B0Y2Hcwu6/e4kgZjt/tPNk+PGmpBCgUP8Mfr+ulS4PzKjvzyRxSOMK6bbAOfJd80djiyYktxvPjt
TfDyEucX70wLFAs7A7CKaMZ+cuTpDYUgXcF5TkHoqr2gn4nfaTjqh7edMXVjWrEJ8co0/A1ySfqx
avbBZcY9z5B4FrldUZFGLsX8yrXI/FSeu22HDQjFiR4CBlAlXZenjrOycXNY+voQMDw3/squsPWS
g55v6XCB+6+HACJpv1GCrp+x45VGlnTPHSMHnu3K+kbkI0ULGxwjR+yp76Xfjfje4f0SSBO2gOKa
IHeqkE3tF+dqZCQfZv4qJlndtLAsyKmfD/owMEVgS2VQcY774Ipb/wXi6IqfiW0LbXrBQtibBcRi
y2rQbhlTGiw98WHrIRzehNoL0PVQbt7pJPREAlnK53BTU7QFJ1f2AjchFTF+d6c+7hK8tZvCpZs5
eYYas+T3AU0QBGgvI+Gkw0KfwFEJ/l/BNOrj2WRb0hqyVbN87LEYVgi+k7ndDUtDvFL5uF+aUNv7
XzWPAGUfCNrOUeTCAjnZAmtLQlJyO0QWERvsUXQteuLqe44whRAMVVCgKCb8fIPdVGqzeEo0kCYY
/VeiM+BYEKVcxgiBkKQ9Uddc3EXVjwvSeLijkgP5tCynRnVNmuSHY/FalGZFcXddpqkC/TudPqzN
2m9sgqLkjrUNjfNnNjjurUGrpDzlRpWeAEEYFfkdkgHTx/X560sanU/E47TnfcndXgTgzbZ5i5jF
TrKgmQefDjH+UvcgLC/tMNDBP3Tv3+xSKGs0UwuIb/bv6nIaS9BVPlsMvmzDah1C/UdOnw8KO78H
fixnl/Apu1ebkWXbwVsnXdywLuQwPPVnHbk28FcB3t46nqCIFJsXZO10ISn54BObpkhMxQQut33T
TF1tIKDl3XwJaN1ALXyLumLLt0WLgwBumfPSmRX5JOQWLfaDCVMXIUUtWnUTyQ6o2DYiW+sAdftV
tbhPdrkMEaiwy+VT8zLd1dyATHRma+v8AhvmCMCavPFMOfrWMfVzdYXbBHzwxqCkb2Eu0NhYZKJS
/7ZNYFxTzHYtoCQlC3wcnM1thk0ybRinvQjQT91hBDldVt+vnaZEjSB8ktTxz01VPryu1/Hi+3ht
pILuyCoxg4fCK05BWZwcSq8+PO6dtloyIXaT4szsR9Wrs2YdRNPgw2dyoYWaJ36JShYkt9ZbCcNN
znz3lhXcWXd8x+hMStJllP0TWKhMnEp7JXxhWSEjSQN7ANfMAh0AstLa5rBC9wBeUsw+CjEgr2Qo
zNEYnlg+r/pQ5BCeAOPCmqKysqMiBr0et6gWA9favjVTu1eEMNEnuLnvwxNQs42Hh3OLITR4niIi
D2Wyda85DjfmqLZCrU8CGA0tZ084c0+H/WKtCVkgUG18eaiZyDbrS6HbnSNZ+6fPKgw56qV2A6oZ
CYKyK2TkypQZ8mFvF99NWnHP+aradkZGLnqQIPTxBvygv0+y37F34k0hTzIZPcltqsslVKEQu9VE
rd9tsvt1v9qIaslfmXrlhln56Q2FTreA5OMwO0vA6yFXaoNVIv7btsHFmdw5GyxcUE2IVw5DmF4B
qnficSLeDvVD2MFthkae3s+J3wOWydATdhHTVV2dxDXLjc13MXIVa+9YFKK8sQwse6+B5tdy2eLP
Kq5Y3Tb0UfjWqobZ8nZ1KiJFmgnbMzBM7bRTfx7j+XsD04MAA8TrcdMWc9IFqEQD7IPVdS+fJH5J
PLPdtU1gGhAXOeSsPHvmV2gkWS+ODr/VhZqoeOHeRZPLTTUoF5kQFKqrGJccVfZn/F2YjUgLKIhN
yFWJuewq5HwBD5DAJcMKD5ys8iNgGyc4MEOFklnvV7jhoXFkm6xuWAkjy1cxf8HG8/x5JXp5b/YB
J9pQpzbDKkn9/s3in4rWqaIXb1zoTknpAhRO7hh2ibxzlMsHhLmVHZGMnS21r8uLOFC4V/e43tLB
Rm7qcfo2tvZapuHDK5xJFC9LTyIKTlRYl9t0SjEnAtUnjIn+2ZH4qnUMFlBDM2kJB8cigjpdGCFR
QE/Wp+UO7PVZbusXlp5LwiokADmcpWYP23AHe8/eFUwziR59GY5m/TuT7WKd1EGJWgDHhvEPq4GW
Js+RyPO+apBYHonf1keanuVrM+hXfUZghKNYVxukVmS2h0lcsVsCsjToEQXAPX/Ad7QyIi+1FG1n
kMeKJvAfOPOXDK4wldWzjNofuNhuTQlVHo6NNOKIlHrIgslYlURCQzUiDjcvMhI2lIv8PkYEsqXG
19ChKcmoGhfjkFwrMHFKzpU75wtnDFqv8hN1zSvF9RVoSwu4B5anniHf8GhhCElb/TgwzZ8fOtCf
bzhL2Ig6Xdun0WqCkA8XIPsb+1j7DpCJWelMpDe78071sNXrxMrSnF7rWvkPEMhLO3lZ7TtIy3CA
56NlECV03tB1xtVtFuMfYJZ0tqZ5Y+jlr+vaeYoXcagXA3CuSnUSbg50D1ckiFkRa2g3iCMjEHf+
3dQyeFJSXyj9rmc4gy3lkgtInWTo9i8JfumJTAK/sJHmD8p/viK7TaHY2l8Su1jA4cBML5bp0ekB
6XAvlT6/sgcGu5g0C7ofT7QlDA32nzAyBAGl3K0yRe4eq9ABHJT3qtfayL/mTRnu5y+OsE5Cztw0
O4/87ulkyIejiBL5SM6PmIU0NLbe1OJ0C1crts6rUHNUj5lXyExo3WYKZ9eynvSxHz5ubkxPoaFh
muWgV+p2fz/OjGpXpGBhKFUt3oKH3L6dqct1oqxmA2zwL/+mFMmHPiWwio1ARYDam2Sc2tck4LoV
/UOj23ORmDqoZQh4JLlmezumLxDTWKnI0LTCZfi4gcMOSrC/HMRtWzM6lx9Hvz9lRZ3uNRXY95F3
i+9Y5o2XktgiJGnYat6cQOyDWDpjxl77Ow74yTtOQzpxfXUX8CncQ8c7u/UmYVCPbiuBsxs82scu
MwBPHCpTiKJDurx6E577mJHeAshPkPbrqAE0bxHdoqHBmb/spC84fI2Y+gLMYJCSD/bL4LxFOI/v
eY1bBaYL2wr42JhWD1HSMZHEEc5BBk/gYc4QqeybvWKNMF8XyPz6c3qoWU952UVhBG6M+jXgKrey
f/IKlaXrFBmsLYxmakejBChgT6BHgZi1IaLM9/O8hDzcbkUcmA6kUcYKvA1XlsImDElPU7vfDl9N
9WypNgE8aO3+pd8q0KEN0SSDNlZHuNEUk8l+SLkJCwMBKZsCfVKbqMo7+MhhuJnNIG1d2CGe55xy
xs770Xup1UesYZ0wuX2kMFD9iJaa1hpzT8vtWu0ieCrVxYfKEodCne22i9tw5UiqlfWUVZraTMWs
tbf4TrrcQArMhXbfUsq4/bzJzDlwPyOsHwRgccXFYcOwFAhHS9uiHFZ6UWqAYJqr6C+/DXN72yAB
09IANMgAGcUed/QVWbV05UxxvPxPxHdfjyqXa/+2CoUGlGQG3JG6IJhj9PhuyUmlQ/ZfeQI4JAcD
j7GWCyxm2Zo2Xof5EjF4NYkbQwILrW9Ssv0xjUf2v1rhJhqbqFiRhxBinG2WUdIE+0/pUGhXpKCj
oDgOBKjRhgzrWkmEZ1hVlILnCKIQRYb4I2J4LP0b5RffzAZFc3XHzfJrc4s7Fq2L5N9Px+ul47U3
MksGgmsTDw075vb1PX4u9hVxZ0rKvTJEBRjPbiXabGMXh2AR4+dfSjcNkVmQwQEtlNOQ6+K6clOL
eLJj85Gy3z/Wx8PN/EIewHdSamg87+s57lQhkHLBc+n1qtrY92Ij2eL16O2S5Y5YaTO4QdREwe2s
CUzUhPQ6X61OoUkLBOFYXegffLqV4HYVLw46MEviGn/wD4qpftSiixKzp6SBIIDOTMa+1Cy5PE9m
PqLvK8HucVRJCjzuY8dsy1ReEUFSvSJdLNGAamMHAx9xayiEopuMS6/u6XeYoWh98acVJ1qF823n
VoTN/9kqnlXkF2C6Pop6BEleAvDmqokIlCS5weRROdH5UN6Ko6NmggvxEgS92p1LGnVuEGk10fyw
uyMFPN5CAinO4v8geaTRM3B0E3lMpcvJImhuTsM30C9wiVmECRCYGPuChonXXpUNYwRQAq2gz1BH
QI1ZKiWG25fjgV9iUmmk8xkH/csp/aGV2+B2gk79lLw5/yXKJXDnOu363PB5GdbA0Ysw7UvPOOZq
/LfjLIXGadSVqxzu8wYEIFae2RY+MUDU7pIYTmLKYQakuQhrhALsmDIMdeoxSeOKTwxOgKnBSxk6
UpiJUoKTYrdj0M0fvexIBTXIQ92CWkq06XcmDdF0DdCFO6Ns46B9BlXFhaLq9Gjgfu+djOi/5TYZ
HbcIlfRrO2+O8e5c0B4KTZUtB+BjzhywPeoWuoVPcazMXjYkmwDWLFHcUG4PooeMJS0S6/cz6L1l
n6V5S9wKEwovi//oPacEzIqLHntWhAzBdm6JmqQeSSDqv9KB0zmWF6/+58Di2PuLVbX/0V91LIPf
lRkw3KCFveVBYLit6wblCqn/TUa4x8zxjRjuG9OdLt6OGuome6SzIB9DXMxHusz1mvaWsObLCON0
zVBcBTeiMfYZGLvN98HBkDerrLud8qKKqZhbQS22eZSKEcDi/0SNjCHv7QjEx78qxA/qX6E0OWO3
FOmYqHW6Xv3CbWMRGhhnIG4wgZfardbojaSkMTO+blfaQhxYGNZf8LxHgRRexWNfU1Md/IFr3NFs
nVrn6TZIFpBHIYYiLNNOOib6NPWrndptugHi1bEUqXqltpXjPxKSqBvDOQS0FXhGLStl0y8uQtwP
jKr6xhqBqwWL54J+SgDqelVMLWCAg4SCG7I0JksgfOaVeQOoGIdgwNieWCd1Y9AAHD8UdrLRKf20
oigHMbdgymZ8QtaKuRG9WuB2irRfHML9OgugpHK0JPywzcDZSNJWBQF6JKfWbjiKt/+xt0YIcQ8B
S2fAvplrJJVE3wgI7CRi90z+W24u8o9NRJJnNe82p42FU+VIMFMQu5d+gr69soCKc7mJAbS166CM
L7oLC3ZXFW3GSEiH5lPu6C9vHqgDL4NAcFK34Xoc8yJXdmxcSenmKLTXKjDzyJTHVcEi/xJ0wKy9
Sw3PdRPEdoX95yuK/2WNeuVYV/zq6ZI3O5E8y/SscTvCbLbncZ9bXEHik5S3+fB6neZ4L+7BeiEn
ssbULi2sfBMl7JUAhrav36VuBPkNgufzwqUXj5zoG/DIyfxrJmRuf9uqUxJIcXjg1zJsjItFAM1U
vhRnh2qSrJpn/BpHrHosoN7O+GZi+R9E1wL7V0grxB83RX/C/hG4GWiZbVvsrppjYULRnaLuyZPi
pxL56Xgep1Nhesjiav38K7iT9F14O3HiJTY/KBAMKbLt3ERIi9QDrvy1WVZEIvn7KBeI8znJjzol
Q5MifpyI7YDifyZwXKoI1g2/7CCIxoAdTRU8+NFnIQPc1NvtugP10verB1/PLUlEseQMDg5jk7Hn
ueNLrj91Jzjp/lD86eBK/Sekgzc8pp6LC8DdBbJZq2Nd2HooACeehzgqNXKlon8TPG5pYwr4je2L
gILxPWMpLeMVrd9x60WeysLLYjp5RqMTOQpMGIifLVv2RRrGLx1ee/aSUQheT0qQiqxZfpIr7FBF
3UKO14DooG8lhDNzoyZ6HrPEbZOF84CvP1AfwpW7tpKP5/eF/uq4zSMRwPvl+ljDaNOYDankIBIp
ByFsVFZlZrlO9jajUs3seq58iqcY21wGVpbi4nRoUKcKrzS2TWUE7Ey/ggTU6avUVk/H55Z/P4dB
rUy0PPSXp7eB2olW1mWJZ9D3ahCdjXg4g0U86fVE1vhmH5RwK/7fh+MGGbb66BjPPB0gfxF8Y4Nb
l8k/VxO1GJhM8VbuTZdUnfMBwqQJa5rac45WKs/X15YV01AEwCiAl11iIBAvOQeKdncEhFH8cqKx
jrr5492MgEt+SUWIYtLHV4Nd0bb6j15iA7AXjbVyk9+byoLgjI/R1wMBMiTUiUJPCYlmciKLAE85
R6yTv36Qtzg9SBz1dLB5i7uhXJdH2Ny9U4JFXN1+6GGLUClfWD/Qt5y7j5XOxmS/XANktMBZ/xdc
L361GfM6Fe2XadKmnEhXznBqTtlKR1zVRIaJ+DuXOt+OoEy5VQ0f5zSFwNa3fcIx9dyMgzJjp2ZE
NnEWvbA5kMQUKANfgZz1sKRqhtRf3gP9bSn77616zaZzISRR2NtLQ7sNru/7/KeJloQuauZ5Ly1k
zmoatTTtIHgUFaXwGNHWUxgrPSVwXjsI2Pcpnzocj6TzYAbAE0BzqTC/mEAy/xqR55QgxY6gr71E
K7CYSjsk6Ul9dsTpxZXqHFJVRpOtzNtP/EOfCckZpnhuu4MapuvCMTFjE1OSxkDEdRFiwsAc1I+/
a9UVE6adg1t79CTuhqjyZvWOh8+/y+elKb5Vd3JYtlRsGmQCs7ED+MP2vfi1ExuI8nXNkKggYamP
HcUxJ5RzBBfv0xZ5M0QMOrWGL66Vspsqt3d9yy1mzkPTtuGaww7cLtORxwpXliRut28Vmfr3AWdi
abeRn0khQ7rLKF9Fa0gdiltHMo/5yE1qfn3IpWR/+OaPn9cKTYfOHzhyqEinfj/RMtYwv+0jr7/f
v50Sg41+001wUSnmwp30+OSJvw+FgW7MsA9GMo0xSeIwyli1gq12iRdrlPwXJ8or5S3G711/A9ea
hukaFvrxR6wmv06aHAAwvyl0aDDNrcvq6kxxFgoXs+wLcPQYDNQXUPr5gbE4jOOR7TwzPXyBgNxi
QiqXqmHHGRHmwCLJgEZ/RpBlLDaoDOhrkeL4MXBY7EfpR+1aWwzp6yxC9rStIDRQScsAucCzV1Kd
Gj7CURh3gC4DI9aGdQ7X7GK8vxXfvM/7B+LCCyi58FDbJ3pkz+8wZVLVzEIS9Xas25wYHjBcjpeb
P2dp7VKuJTfokbGfsqQKSte8cUYCBpnrOrl6E3LHanrthhUcTB2pXO2oCs29wlKL5MwA6Ptv8+OX
O0rKeZzFEXpJOqmE2eoT+os88dW4EoTcJjtQ2M5Btm66ghVGWq67bFlh3+kFyoMVDpKbugd26Wdx
hwNMqcd32WFzkzHd8SaC6BzAaNX5GcBsq6L2+27Wou7nKiXgKkUvTAWPJseoEgbNC//tWKmkarI+
ATzTLHWi1kWclmJjJ5vHi2/OIUouj6Nz0k8JaesBzjuPQfu+fRoto0/L2w+NglCjELk25doaUbZd
fMDtMUTxoFCGfg2GX0AY345+C1+D8K4L8EEfVl/DQougeccIYnEpV/14alz437ez+budh4lGGAiJ
HpwM+KVvjMZ/WawGhhXzPnQH9kQjdzqQiKw9+re4DewHiDmrVu8DxQaQMHM1CjfHpp1XdFvtEhT3
MxeCnFMrnHcgtTtTLZRHqPj0hDQJEF8V85bL5VKqpHWoN8pcT8hz9TBWHUKrUWlTTfRviy6epXEB
C2f9pe3QMs2uMFYepUMnw4Epi71XOoDBhC9b6+DpPhsoWLBOlEHH8S2StDhj1NFv0dxcem0rjhmm
IkSsD6KsW1RKfEo8d/qrDTNn59asy0+qWUpp/Voti8tbRr0DOHZGNoY/BuzVc5puWgKGnl8YSg73
HhmiUX7AzvzzJ0fKunZPr7+N1AAOp+hyFOPLNq2IZlFbjrA9M36NJHj9ZeJAWpotu4XgtDcB87QT
DZMNSEi75WlP0+OoYHZsM9G/FkiRz+QP0VYN669hXLCXInqCPk8fDnasDICyRjWro9r+zuuQLinj
hJOsGfjtcsP9uE1YL6Ev0aOb5DdnUk6NY6ohuruORl7xt7/+0JEyioD70Ot0aiACh1xFzhR18hNo
cfIoLe7Ew4wyO4+RWlcfyYzFd3iSYQXPFne8OyuqC2iZ6E3XYXMBVj6GgpVVi3Mu2HfSGS/H1JuY
IKaKb4BilQHOyuThXPHSWAggU+IfcFL2XQDlUv1qclM59wrRlRJ34LyBw3a14PODwu15M+kItox4
/9myxa74bXNwZ9gy0Ms5am7Ww/sTJvnjg0n5k89Br93tQSrjgVj420qwbaRFk9g/Uxg/15Uqziki
6BAqnlnlk7vdT6enGkGpiVR8bfLsaIFI56q6MQ7Dnrgqmxxhv47Xp1gbiFAL+e7kQzHroD+TvfwX
bSYa55gID5a6AiBYo34VZkEh5lZdIPh9qnnp0CEIAlsD/vSmSUhOss6I1sJ1rrc2h/joVUcNrMlH
Ha/8+ou+a94e/sS6+kIYo0FY7JwCu3DjSOAjcqE3Z3zyYGa1pSlr46PcVL6AxYhy9XI8yJ2MKS0Z
7GqfuB6Vcv8p/fVIj/aj9WvxPGxyTQR3J+ulrFvBLAmoISS+4AfY/0X6345w1BUkpOkAOjvko7s5
4M4QcRIn4mYV8wgIBiJ27a2Ta6Bp2J+NCWRlpsBB7T6RIvkQy9+XyRagWuiKxL3Ff7TnNuXs3S9O
DuKHcjdtJvTNOry2SmTALJAyBuQkgq940vHs2gdJF9mQxTZ9+FnivM282CKYrx8+3H4E5VIBDcaV
VN5pV0t1I/DLtrzbJs6Emn7cywbU+Rewl4VLjDBgKMtZwLyVBxrCXxGHy2azGMac1XH91w2jfQI4
NH9H8Hr/o6huvsFPkN/kfiP8qVOHQSWbuCpQfh48vtd1mdLzujtsBBuBLlk3zN7bzpicBCWJiLry
oeDBl39dcNW7/v6xfF6IR7t1riOHl8MEkTjS6JIH+vFnDVFvMWcYxOegppDctia8+hSuc0i3nLCV
uPd/E66RNDqJyhayiaDjvIoTxD7zOnjx0yq6DeF3QVNZyq0hi5AJmmDx0JkOqgH0uhB6tdJPmgVZ
vE1yXj755j2ds1Ii8HyBPQK0MLlOTCBNPC8a2RIvixjQltVV37KIdXHGJvZCGJCC2ZXSLsWzEPbC
1Tm2zrA30dXrnUc4h59AiUc25H5XZzCxuI2hmC69VRNr0tyVr6gBR+qHFrhq0kKuZ81zV5lB+hUn
5u6/D+BlJzfY+uvHDKAC3RpkNF9la343up6JSsqlsPSGOI4V7wQh5OvaxaxeCNfLmheRl26LZ29i
8RDZJEiPOkKZGGj17a0Q3f3GKzCjvVMnAnzJ2r0d4umAwpXZkOCHPAguFVWA6VLy0A0dLEhv3ZiT
H4SOd5hmVEUbAQGruK+FrbqX6NZvwJGPCMj7KNpMivihK0yQUalE8b7NhAbIBcumqhl5Twi8Pnpa
rMgBpipAmwMd3TClOgV4olXvGL/KMxP2PUT8FFcnN+iy/uCyj5rav1wabQYCVrKhReQwixQvlQsw
fpExExiPWjx6yXkMtXHdf7vHzz28ssRHrNoJgsH1Ytt6E4UQNXb0qYzFYJOnae4Am95rQLh2+8P4
AZdT9jIoqGv5hiI4YbUcX0QD20Jd7f5Vy82197hlqg+pgxpxsxWy3cBoORdBRUciJzhUHRGHr9CI
905ZwNIbgBmMqmc/19/uJuKUcTvJiCup4qbo0PIsNVAvIGpGeJyUatwExiCOqqeZMGzM3PUMZ56L
MM9jcUG+oYprHE4MuUTZ4sN2ux1DPD7JAAxBNrKku5mZWlPmyQkwz/dXjEG2FERLcxjOlc4IP79s
d40NZ64GmrqlRKxpnkKQ06qOA+WsbZhmZaKsKjWeI9X+sTHiO/5COVKAy3Fzu8jStJc+y07JjSOL
nsbpDZjLjdG7BRZckcOtwHKZadlGYG70mWwttEcP3RnL2+0RkPfha8vdwftDz4IYR2a71pFBDggZ
nOcp/3Tj9yWRUbjIdk/YC7AKCSDp1rSCQqJ64OYlcLz5fyvwBhnV2Q3yJAe6HUg88QHlb57ctbtf
+vpXqgWw90qBkmhn2jF0vDg+F/2wJl7ItMpTehHCH8r+tMRMX2+Cj0U3eujAJ3BoWbzMTOgw/Gks
TdKk33dILqaSNy7N9FjHopIAS/uteZu91Xk3MSzCAA26vVUCgpwPG4S5wyx4lqemDj/vEs35ViNz
5XODY7mHtvHgmvPnCftLDwPm+3Uucv9bhL7g4/NtxBMX4iQLUbdXR7zsAJ6coy7MTNYjfv+fsaYQ
nNSQ/mhivkIVsypBsrp0QpUzNn9aErOR2Jooh0RTJPafooh/863DhHnLvFrnUAiuTF4/XwVS2t/A
PvuTsqjCrI0/oyzzCo/mvnl+5qzurLeBBHlM7btX+GIQA/NLqrPakEHdTimcdi6nM3pD19ubWjMW
G0eI2cSKWqTH1PDoO9laM4CakFhbV7hPPXh5FLXn9UoaiLJ2htuRegjZY4GbYX9gRTWedQNfspnW
lw8bR7jIRET0xl4RR8itIIpMg1hUyTZKkKKXEFfVNbDqv+OaUg4Ha68HDjHLF4RdsMCqOZACdlVs
4i6pZkDFOpx2rcL05SvSmy0Fix37X8QYHL7z/I65K5wES0F4wIuWXns1UWVAx6a55QqqG8M9jrr6
CDl1smpByprxjC6yhRzyreFTuU9J1THVr1kA48/psi0ta5hA6k/aGPxC3mLNdpbrnwGG9s7KF3ZA
P68kmGehJq0bn2w+oA4g67j0/252AP/TEPxmAsL7AjY6ZdTSJn5OjBgxLYMOuMxwaVUKX3eTKkPR
K0jknZ9dm0u6ZHR/XqeWxwXwCjrR9ia9/Iq+Sv/4xJDffWhlHfPT9aBj6Ukjz0rr4CspH2JyjGqm
B4CGQJn+vFV/njEPxCeBX9LmJ0MtbM7BnKDIUFQG7pK+ORREEc60rnMcmiExVfAyTQvC65OkoLhu
7tfiwhE/DDCo0whlVQczgfIDzaNumpNEtkPXL7wRMuAXJj/f246ndzwP1MxZhbXGy1lDiuRCRgsm
maoX1upFviSuE9DlSih3moxeE/HnE0FYJEAw8MrsKd4O5GGbjfRwfU1BtKXeqTk57BhN+MozNZjP
piRKKfCDIoUdRs6Zf6MR3zpj/rthOY/ZPYvG0mudBbpvVOo3JWsjzIc0JR6Z/VdpVZ1G31PkK4ZX
ZhAXPiS0BUTH617MdkeBi6YfkLwe8CzFYNl5BWpqaM1u7ABPq3wLG+qbJOx1pqXookXEahkdj5ZV
q04PGivEAfMwgFnJDsh57jb7BDe9nMkpC9RgvKVqLMEjRW4/Jz1omy+avt2GOY8pJtG3Fy26RHwz
sdvofMyYLLCDLhhu/vRDZf1kLgXiujBPdWBO3EtFiPMghEHf5X8i99QsvH+Z/LcWfwaNhI2ncoLi
LgL6nshhkJk7fmHwiK/iYpGcpEnmgS/eMHmGKwfSNE8+2Gm7ldKvP7pESFLsnbHN4T2gmMh6mKzR
SN8RCCQTnbM5JAtQHNR0zorr+Glx2+5UMHU6jmVwoW7ZakgmoGPh46P6nA7cdWraUoZbZBxCmijn
nwcVHUS3CtijlyenRoZAZxpSByXaEd60cs9j4Fr3cXEW/7A3KAytbE6/umtPgkrS6bkGvcLx1U2b
iroxvia0qpipDKHOjq7ey8r9pKPwzh5tcysvZPQn0xHrbg+1jUWXndztsyFXu2Ktgf5zWz6k6CQw
wZM7ykq70JbohCae2x86eTJ5HG2RhlcTcCUBOQLIpLY7c5n7M8WvcicLcfQDzo2UUN46QIhsVYKo
n9YcxDj2Y5HPsBDms3rXckwk48aXMy3rUFalcpdaRyRQiOWGXzm6jA+s3BWHsDL98wbrOneM1uBm
y3nmPNx1mHSiUVl7GvkRqy5OGs67VsjM0XKdd9hcBz7kYpXspOmAdjHezJvzrx0qDar2HLTlCn40
F/B+rv+K1AJtSsw4J6PTEayjCCO6+5pQ0fD5P0ifZMSJXYY69QW2ycPXtIgfizX+C+5U6Ctp5B2B
wGIfcyJlNcM8AS6nUYs0/wZIDS5kqGQa2uZzpN1U7OusRC9XjXMNFhTS0gva+mODTkHPwKfNSjrA
Y4S00iEKnj+Q436sQBRVqUNqMnGBZ66e2dot4eMaVqXkH8Dsq5gE5SI+9HTZNakVDcYmOpd8UCli
nIggGzmN4i4Cru6J5ioRSPDOI3uv3VBIQBntvN6z/J/QOIata0ke8T1eu19IipUSD5O7IU8JNuae
XXGlzM0aRp/AwatLXyMRk9pOkAHmg5GH/MMyL3KrtGXTW02qRg4KD5vtnPBd3RAEfc1GIyOF2Ok5
qlhxgevIUkU+BhW6D3Iejx1BYJ18KpL7Mn2dz4jMSWs0NdnyRM/xHRZgGtDMBDwl0E8208xP59XR
uPh/No1mX+H/y3/4V9ArUNL4oD9g06gyawgAt14TqMqQQHhv2FMtpGt/TbCL6cCTf1KdeXKHv260
TiO1+B2PCXG4rLB8ReVveFrh1CLgk0VnHDOrQ8vUq/2UaIJ70D6YDq42v17wmySv1cPT+44JYylA
Q4TWtespldkD7wfO3NlQNDIS7ArIE5s5PSZoPIfHAf7TLfSab6mDlbx7n1e6OEbVnW9iMbwsqQJC
bX9o1OHQ6ajM2hVlwkq28CG1y6d+Fm0l1bMRDDOr6mNHxxEXEWpIqKRbXQnEYbdYY8pJBy3fUvFM
1foWWPckxh9Hu1K+Bbyv1I9Mjg/mTMkiOqgLNNPcKAMSoulEof+nB4AXQoHzFlDXxaOorkfVZBp7
oDiFBT+GBToHDShqU7wqCEYMLh1v7qqC2so5oc2fCfyrFcRZh8CdxkRfjHLWofUg3nd6AiQ0MoER
GaF825ecuOtgB4glp/MDcBrstOJeR4toRWqu6lRNLJ2IFW/H2fysvd1R93/WLvG5/dxzl6da2hDQ
p/ICfbxy3JWurDneS6XZ6mQD7CJDbX9dDVx7ryzh5G8dRf618rluLoWMeKt/YQcZmV9Y99pmuTZj
xeWMavgUZkMC2Ilc76d3T4CVuhpgqd7Kp7aCay5DkIUHDTImDcq8CqvnBJkta2/SwjNRXtvPiZB2
gZ3u+uM9tybbIhWOtYmYTqJMbUgYNLNBfybi6Ong0ZKskBH7m59OqIbmYCpXQdnIOhp/xloou2V0
uk1K1Cs3ijPAJHI7gXuZAiSlHv0ge1pIP8m5rjyTizrPAHTw/5gpksy3U5cqLnTSHByPnkqC8zUr
UB4EJpQImbptv8kkuN586avT4Z+EqLxJmtG08JFl2QjmZe9LJgl3LAMI9ZtCSx68f0L+9QJg7jWK
S+2LoNhJhq8vb3R3OOuAXkkfyxFXNifZl3qm2SRm5RpLfplWhtXN/YymEMA6z0PPGLqvvYNHt8DJ
vsGfSCi3QQbjX/olC/Z3SDHeKdEQXakRsCK71A1NTkjHJ0aeVjDX6BgfTa4kcK0nxGZtZLrL2ZUQ
ejdxuOBXJGWDNIOe4Hcklny9WvoTMcz6O1YW+EI/Wv04g9ZMhBkIicJPdIMM9cc7k5LvVWQQIvkI
kVpuyc4YdolEaNIeq4sNJlNRiZyM3bmO98z9aqeH65U3fVblrxolHBSfBmk6PB5/Qk6gVnLbZfGU
JrApl60xYDeyf2HiMkVoy5V/NzNfGMtl12OATT4o+utVOvAKc/kgy9DMYsHjGy5yvLU0MNYqW695
a4p2ixm6QDA+bclu7PgqiWbHmbM3iygPnd0BFdWFe6RPkx3Ysh4hmcbvvvIHFjDarqx9Y2hGv6ho
n5ZGn3At5Wtg6SwnK8a9ZMhMsRIO5KwHTZgmqV8CWquYXfPz3aBWzJQAEfABo6nX7N8OQlB6FTq/
XF82lecH7od0YUu61N8r+trFlRnDXm2s5VO4kne7Lt9T6I6C2fVCODzczoiT9b4WtTnelsYPO0tY
9ct/St8tHapDNNNKiOwcx0szHEcthNnjBL3xZEGKyxD7nm92tqZeQp/BMiMB/7uu6ql+GtOe0o+X
/0HZ3k4PNugkFoadIyI94WKlh4cV08xiHiZ/bc9YvJ+2AIxSqsTXH+OclblBRHEnu+Mec3wqqgKK
2hT1TnEiedaoLQyVWnoDaASGRQS7trOCrxeR+6rpfKFBieTWGrd6oRr9lv7fWBdizCLg27mTPKon
/muggu9nicXxOW9SpuU4o5Oi2bniC9F2MnueC/Y26yAkLUqBFNiq3aeemCeHQudYdVfynHoL9lbe
MwqzXtpxampXeCwZ9o4hCRizJUgsQJQEMwGpTaGNvC7fb+RNwTPSBnRRtZCtlGaiV8O5MfVm2pT4
nslkCahvpYhuu7AnTqCEfPmhYJIRwhDnfqof4hSQ4NHvXDYbcTrFRcD4v04AOpPzCbMr1SfPOtS0
N87ZL3SCTqN4LLoEGNygPvkoRR8JXpQ2jFyXlQTj4rAw3AO1eF882llAw+FzETOoFlHGfL47QQqG
lChAoCwFJ9O801hsgAG1fSv7owE4QDbOHH8/PjQA3+gSE1XC9sN1fqTVrYd++k5YwE6yNn82+qr5
idz5PNstblJNgJBcVU9/20kw0eGYZCqDkTnxJT5ysHSLBNKK0pid81SERPE0waexWiQxeUewlMzF
X8BCJe7DumIpLdGCD6sStfbLTAVT7JW0AU7toNT0wp8w5LZD76Htra4rTowjVKpqAYl5Re0POOQT
exe34pTFbvZvrCq6gkBruqKE0GfKL1E6Gun6o/r7BKbLazgUbpKeby9IqXaepwWL/1Ih+qMjSvMb
iU5og8kDADjjW0JXGd1DLcFO26h9A/ZPY3iutkurbw82aok2gzaNGGKwglfjAXO4g/MjdhSevNCP
jm7o3BNhO0V9FJ+xyxt7pV/r8R++DyS6LfEh4TFr7dY8Lwc5ChailWL3RGiw8+PHq1aqZNuwxrZ9
1WP49IppCbgDayWizpzFAFHacl9aTijjAgisro/mqW+8Ec1GcW0tZQbHwMnnbIo3YN30fNLPjWgA
TKVxvIoatF2ex+CQoJ0C6jVU2cTRuHZrysy7yT39vGb6lhgHDVQAr9r74qDkgQkzg3fXrJ2F6oyX
cLCa4RqX8Ckuh19pjU3zXh9PcRXtYmEkEcRXZWSeOkYc0k8Dz3EvW1oIRmdswv+N9hGglE20ahbl
cMOsH6prZatV0Ikry2dq+96ab19RMrQWLMUs5MfkNVKyn/MxndNUF/ECD3gRBjoynjavVZo92eHb
YJDVPeYDU0bVwczgWx5SsldEchiXEu9XUXq7RQiL9XLnxBL6bH0e4uFwDEKccfNEhavsvGrsoaPM
w0uc6SB66Ld1D3tHmKKHjeT/esahzvH9ueomhGWAq8HcocVwNx89J93A7EWaVvq8QRLoSOk7rLnb
eFk1gfVOohBsQ4G5PRJ98zsat2dsYCfxcBDUfnp8nIi4+qJmXvTKCmRShwhvTPNJLOI1uyMtj80H
AQreqXG07gr6vSX2FBUZdb7+GkMU/f897TLBNABTzWPWSoeQOLZaFzgrPwOyxzNesfxxDLN1JmvS
9i/3TwgHxV/knZxI/pt5p1L5RG1p2OVAnZbziSw7Aiomd78cuZsoYGqPEusKU44bQxKViiTzKccE
BYUKWKpKJpyuzQTvXw78WqNvzdnF7XQ2dBFguSbDMqgcilxdInqQMACCOZW5A1Y8d5zBlRu1PV4h
lrTOVOw4XxDJLROT2mA9oxcaZFNcb/cHIe4pxWM21NkJZKfwjXckWdEJ1iyl6j1oXHy2P5PMRGLX
kCVQESekbJj9PMUM58t9S9qwdQhQXJfxpKtO3p+/sOek7FOQj3J2cywQ8N1kXuzX2/S7s6ewTLg3
UnP4s/2DHedBDzFNsk3eFHtpcOBj/4G15vBJlbeyyIBFu7oGUY+c5P5KXHDPXn8RkO3IDwhE4LAy
UBzp8a+y2VTcPJ5xThDnOYKot4gIo1YIuAkCNaIeHLsIpTXX4O//LALMoKuGJDyWR8ayqcfZWiWz
LGhKBiDfCNQmSEtvATXCcGRss4ekbkGKAgtrd5XIbfPscx/hpRKynNmGFmi6wpNxwpJTFeTU7oDJ
6/6DZRD/DsZanV4QUjcyOJb14r1ZMdL4bftgsP/OnA5vD61yTiVwzGhzmhSD5iMw05n1ErE8w7hw
ySyjCVPWATSp1aORemvjIhjenwh4RzzHFSZRfX54c+O/Uh10LgIfJlfDvq6SBN6jBhtQJqoP4vaU
6g9++LeelvcYxSCXZ60pNMOJyxXXD8u1LtzmopkyYqChpPPRPa70CWdA47s77QMLsisCYy5w5ezC
grZdBl+k8xu2owg8bh318j4D5C0s/rSoDpwItmkS/KmwP3xvpQJGM+yWmKpNnXYpcZfg4eQsKBCF
v3rGDePTe8lewtvmjCsynJh5BXF/M8unF0T7dmbu+cRHQk+letH0UgS/5n8Irp3KpRUwHcDnhN7r
0VjMW8JTeFYvR98Ajruy0VqSuRka11v7eGHlzwkmHkBfu43Encej8YXFS5QjY3Cn5YZmpgrzZCNw
d9XdI1pRafsvScPFmJYeke/TpnHV4z/wTqmbQ7NdxTIOh2naMcOyLOJi9GZhhxLvIxlEr2pXcgg/
El9wc5ahB07kE81Z6QYA1dFlRKWEODXi6Gp4dTIS+2OKkTbVCrU5bSIHNRMHtt5t6YxdhtbTjtfl
7xRyDVECISpO88TiUPY90YnKL1GnahSi1yfk02KA9P9VNkhC91AL+ny0JHBr+g8oBAIcrWw4zJzT
VbqFHbndG0OsH2KKbKttdShcFyqwEPcI5IuTSPsMQPB+pSV/RHdjadHIE/RMNuUpCaB+H2Bembwa
z6UTm9EGW7dEZclu4YViiy5E9I6Pi6b3+QB0KrPuWoFo+fS9mc9ct0GEGA/vyHO7GwXZjccUwLqb
y6VQZ8ez6DU56yMFXKzhUMjsk6PHya06rhJMDfLOtfTZ9XcKx0GEHuG0jUytddqZKJx3s9tHrwLL
rb8wTqPVrJaZvj5kahS/NK6SF8H1mq0A62R9NFYTcK2v8MSuo7tYwzZHAOMpguBq+2DWLpCiA460
qxtuYA5uB/RrsaBgo0bZbGvImEW6ovjtINcy+bKeMgVvcdtNtpyVnzUQDel6YJePwtR6M2N+YTJw
vROQH+3XDc2XqsIJs7mrHLXpAFKGQXgORoEiWpf65aLEgpRXv/Uw0drGuNoxGKffX6kC8IuNBk2N
BoIPNJiEhgSP7IfaojD97OXs++110zv0elknNe6/6EaSu9KelIkHekU4+4F4aR2nKrt1HnKA1zB9
LGv43oekjfUFSlZMLZHmptagM5bNacZU6BmXyxIF5F3Lb8JnkxUtTFb6kOqSSU4/toI2K624lcEo
aEbbf+1DxURTiA6fMJGp9eHUpMpKQs9p5fHYyvQZE7gQoUqhwK72qkJizQpFmh48lbGGiFJlCI4r
g1Ua1dwHzFmHA1PhOYoeh5iYtq6cDNacJh0NLVXq5rSYi/LfpKX6LfvGSn6uHyXiEnP9O/tUOpO1
JtPcSJbg+BqrOGUeTCCzFB/BeCMYVbOFNccdcwJkjNXCSqYkQtfbvPP9Ei6ou+5Hiip2y4swdaFy
pOrA2ZK+AF31HbsluMYhGSWyNGEyM1KEGk4rVgK3CotxqyjvMNS1cVPquniirAa5YYrmtbyNaUrR
lqJVMDvXeUNsGbuzsaIVYorStGpjiVcdWBIG86vUUPO/WWZNrgye7rhxccAclRpvvZwSnPWRvU/4
iFsEpLuQhVbtdYBxu7nqR0imu/CT+THDAfxeT7MbCWQ/0K1KNs8oGwwobEfwB5V+Le+Mpfv0j8J/
pgWuJ4F105afqJ2DgTE5T1rnxXdjx9XPpm6Avok9hgPbh8yskMCwzv7fGdzgh8cbkvEu945xb4Hg
LiLtyyXiGQspjHGQYoEU7g2aFesItU2y+jE/VtKfp5hMDrm6OL/T1DGLdqQ+eCeDjNrEUigh9u0g
ho5aV5FX6xsBHomkXRS2MrXMwoHVwhkluTyTfwg15G8rDGeXXcw0V95o3UtOuHY60mOcB2J/0KFL
neGBFAsP6ffbPBxKE73WCNL6lidXLHJjYLHZkJp11WPuktQleacVK3VS4DLSEFIyX0/w9gZLdUzF
7Rchx8IGnjhLC4KVqbwKQYNeUWHAyYApZN08DqveR35f6H49B3psjKqmaNezrneyCearKWcTU7Vn
O8HpXqhE1b2MN1m02tf2enw29d2ywtBUY9XJzKM6mfGSXey0q0P6sEu6rT51lTTFthH6geVVSrrK
wktuG2/yHkk4Iv333cq+MuEYjvX93mMMGDXgK9mSnYZR6mk237ovKnF17qN9IILIF1ub3W64zce1
pTZbeH7nmve8eMY1g5b4wHcpzUN0LqYnPxch1XTh8HORO35uIPGLBICvPklBsCeDgBYaaEbPm25K
nIijdam+b1gyziJXp5FrOir/xeBixWjhr5zYHAXjLQhhrqtbmW3vsUxI59z/oq5ePodgxo9JxrIT
0udDKfn7afzQKYRBQK2yao7jUfYPsRHDg7YuV3XzQ98KBuLLXUo7CPvKSv0OrHGyR2guz+omCPLX
0kyxLMvtrizlyuFgn3nZ2AZMZXnDHiUwglLEyo7RVoKTZCxbY5AefBRvHz4OzDvKffjK24ZF7R76
sBjzp7mTzMlkHkm7B8hZsMl2283lhwRqW/0hEpnUSFM88kr4u5/hh15B2mT6UUyguI9Xv1Oy+8no
bfElFIyYaAMGBwEdDgk8aw4s/ZLQDPeUt4MoF1J5TaDSERC5EGtLZ3uGAPAydSm7pfpSvagtp/3b
m6aoCjTZ58gGeSNRW+SEIbUmv9Ggts3y7iBQOSV5ryhJ4qIVZWXQ8lextBpcEHXil55TrkaCUyDa
L1/8uHWr0ii4/M67sJ3RqjqLSUd3JKcxL1Vv6UjjXFEI8QoEZKjrkV04WKHLSABEnNVnB7Q5Su9y
beGZ2+iQj/OApHuowukurUSbo8VlV33ta1L7uMtL2d9Y6gMo2S8fFTbPCW8Vw6sb4++Y2j6gPWhl
fLF93XC3EJ1AyvgdziaJpk4g/QMEGfZfIV8Q7dGUZ59Zmhrpw+FFmNPg8YluPE7I3ij6AKYOkcnJ
qoSKUiPXiDy2ZX4l28rXkZlo/ysYP/Byb2ByvVHia9S7dP0QuuGrAFMP4+9lXO/xzm1ESSLzTQ6y
z7eLHSHBFROYBzPyweB+i9dhFXE7u9gnXBx8+F4A6KLJKcXDoIfeTF0SBn3ELz6/aYvCfz+/YbhV
hpjhszChgL4bpn0JKieEsDFx/x5wbj87G952xmAoVcPhMymgAJnYFre1t7dOl6oKJVAa3gmj/vLh
c6oknIAvkrLu5pzvKJvtyAUCYBl/gBzirV8wvyvDjhJn0l08lK/ELq9wwc/6mqjUECBbQ2MPDNZW
bvIywaFTXuWQW8sYDZCiJl5tLm5HBckOb0aWHNMlkaZOkEllH2kPWMHcwMgZZSRLUcZukr4/sPWL
jdk3lVXYYZu4KoTwc2qa5ANHc1t/UTy023VK/pBzu0t+qAoduq+80v/4kSzDqyvSiqealYmBq52O
jIGppun+WLCQHklvBfkpD2PGCBwrCdPJVWy0Zh1F4UWgXZK7scs3FzLFSNRxHdSKcumL59agSe18
EGxF9d03dFjd+ZmXqxI8E0tXlhUPQUq2Q93VNOJ7x1xIDxlGS2SRFZzzq7TZHqEYckpdPqjAdSTK
5k+JLqUhfv+v328hvp55+421sITAevVpZAkMy7hsceblOlqk+oXoYj/jmEnPGrkmqAW2XFO+oeCd
AHezmd1+U+WcaplA1t2BnUKt5RcAQutSwwp4lXDr6wfTSHcG/TlhuE0JAZl5B7W7miSCbJ2bJIm1
HC9mGbuNgrlqHW2ICuUuAiOSlbP8tc8567Edm0ARPGeqMDHF2++/0GXJPyxhUxQtx3K1H5UjwDBu
qQJQD32nBh1ixhMixmr1o8edviGCd25ltM4B3KoJ5XTuuetKVYghqSn5PraOp5nksm6HaAF/r1iR
Eg4Dz2xCF+CVrJ3imdbC6mDyeZvNhYE+6jA6FJOp63SrC8uIcBddGeE4OTtpHK2Y36mtQn8zaDdc
nXpto61e8Op2uV4auLElcx6gNa5if9q/+ztcJiSE/mC7zChyCRyGNGlh/2xKoKfCo0B7MXzanbRj
55p1Zu3X5/BWaVj4SgW58isNWUvh7fheJW85BfETh6k3+EbCDw9MkIRRqYNT3JWPh/yhoJce3qNz
ZrOsZ9Y+n26z1kJaZ6OHxSNLQpLKZBdfJ7e43uJ2w6mom/dspywwHXFa8mEBf74wbBgGDWVgHGpA
JwJ5bL+MLHLnXDzoDfcDm4Di5EEr/55scz/5YMazLG5pO92ZJlxnzmu5FAHiW3K9q44uAeLdlJyD
jSQvPEXeJv3o5nyFBxCUwKFeGlQmBEe7T7sGYgL4v90Guk7/ZphJprodETEWZHAEnlS+6hSfYkDv
hgKxQzKvpUGEQSUT2jAmezyX35vP1OmtU0oeXW7g4zDWjAnye4DNSsHM68vsn5vSjyPqeewXyNux
dR6hGyJh6fLBkRUh9NRMztnI7r19AyOZFhTA5LHu3flrzjhqyj+Joq2cfA31yb4yX1LJCwJ0F7Xa
EPgfw+nCeEASPNE3IMw0zOoqhzAq5SoqnLs3HLqNyXxH4ylFCJaMlbSUM1r61Er/XegF4XRJXxX9
++C+CwarJC4Yf6vOaGUe7hUMyySM8WaGnbbVdH3PaCCxk6DdAHqGd8aMixhR3itoHFlRbxwSFEgk
TdE7zgLxh4x9PfJ4l8CmRNHeiMVzlLKBdTLyQuJGEdpMGDIL8HeaDuRJntHD42Jr8tiL7eyDzSq9
Gdcz88TsJIWa86Yde1liUpmUlRuPs+I7PQl9UYvubyVD+E4HD4KWQkUtpY3BpFXCZ8op97lmShmc
eCuOvB/A724797PdAXkUdh/xDXkP0rtkqdTofnP59o5q+5nISEGpRWFZ4E3SukIHANb4s6pqGYQu
dIbztJRHZDd4WED1buc7og3vhZFDDAWeShNN/nJN2xHgqKl3YNfNfH5UXoZ1Mj2OwY/TACwNXzLd
O7vZU28cRpJPJ/CXjp/t2qOLNSv+eMTd5QTqKW4d6MAsx9NbURHUcvUpXKio0Zi1hJ/O/ftPdx5l
HSNw4rAQq5oO0m/dFn6i8Z6lfGInp+JdJS5FDAuiDO6ZOiprlh8o2FMNRmlPz7ggTLkQ7W2rFnLx
2RI0mipIH+ff2PHuh/rCE98xmtS7ro8EO6ABkbXbVbJ1qw0/cYo3hnS0sTdtXGgvPDtaihHN+q1T
3fpW1pLnhRNHaOfy3eQQaz8KHOal2IOvkAL6lq6DYGYmXFiKCUnDZOzeSBPSeYYeeASXC8tDy7OU
YbCAB4tmuXuhbMQWVQSu6jBq+q2eiM0J5V9P2YVPWQx9OhZF0ppwMAsXMnESkmZSjkBwS9F+1o5m
+g1VK7jQJEC6G34Z3EEIYXr25xSrViMF/QGdc7ZXcz8y7NnRElCX/rpmo9GVuqSu6aTm34d6C62n
HXP8iHA3gi91IadJYrXuuDdA8NTPT+i+12sROnPyBqoqla/Uuis4RrAVsXsqNMpM+g1waPXSHWhP
cSsf4HTugjV9RHfqbQnBCgmHqqFeERw9UuWZXVXk2rdGspSGU/1zkuRUvWwNpCZ0AkLhWq/3Kwo2
xy42eicp9i/QxrkK8rkjj2nU+Q0zDy60Tb+7dkhD3EiUgvRAUx0B8z100wMN7Dz2GUziC8TdVll4
1jV54CrHTpV15iZUjUV84cn4516v8ZtT0iu/psP0oHioomLbu4wLAmwDf+B5a4eeDl4dyVIbFcrt
r7lJtaQfAGDPBcUcWaUIXtny5reo0grFDiN633tBQhxx1hJ7kfNWJsemM2TaUMMuxdeRH4ihgd4r
LHCx+O6UwWZCfBnydwMT4IZvTN2Ut8ONYEzTFm1pW2D63u1h74RaLGgOIj2nQUfMkK064gJLdhkF
ydmz/h+oe2JXOKvxMNkTd1OOf0jbQl8IjKb0iIX9mCdeIyGWiQiw3x4nULoJUm3MKZUyvfnOIv0M
it+X2UJGpG/CsgIGZa64hlfmyls4ghsGhhZZxkWU2Tfk75ZF/qUKBX4JhVXRyNc5njylsdO/ieaN
S+smVX7X5A8r+QrLhX4/nEyh4b3DYNw4l87NDqH3cEeR68vrEKAg5r5yAlDvqFxasYRFjc8ZtO7Y
UQoFV4ifPNH+2O/bsQX1ond6GmKOQLhDT63YdcfUAyeN+IP0UgriyN0HbaOoJchWuQ4lLQRqK7Qg
Nlnt71QtGKZ9sTIb8Ulh8eLs9tdYts6IJCxP8moI2L4HALucIgegaTzGG5TITfp0yquM0sMa/yAy
uSo9GQZGF078+udbhCK+iO/+BIQwvENRytagTDAFwhG7tNK9B123ljO+r/yyR3zm8oW/3AsqWnKI
9Gx/iowqAPCu870AAz+LLL+kUUaNpRk6V4v7LC3xQpc9CBEv2AXBISYrB0HlLP66rfM+YLultb6O
rsn7OIFKmjXy5cxgHY8lpGgfUpsKwHl3eQWj8PArfMbhY5PZGX0iotZR8wMScyGy+RY5d7uD2pxU
0NHZWinh7JjKgn2Ae8xqDLre9vYuToTE1tbfTq5QVak3LQMHSjlifzpHFR/Y/+l1s7N7gtpHoPjp
dT49Qapu7G+KsX5BjK4NQA8gQ7CG4pETadUnjvuA9ZW9kMqOWyKp8BqfXuAYAk6TPY+PKN+uNSDG
r/oCqON6wB/RSTdKzZStqxfFlQV33Z1fbBJsuT/S82sMDWTxf9mrxooWL4Whz1DTbpKPdAiJkygT
rd170Aa1jUVXpMPtWCWf5NwSnRNF3sjjA0HQZib3m4AIOcayoPdlcG6ydbtGkwCqsC8YOai53eun
ZgNjWfIc3hP/zjysCoDFYnN7Ft/KPVljnFLICHPzpLLC1k8A1e9jS9YWHS1F1jqJ68BMyy6POzpI
qB+rIcoFDs2OXIMLAUfCbydBiMddfzMMa6wGpIvUakLasr7ddphBsRyFndpufohVemsaBDsUeEn1
2dtjUA8hWRHKAEbPR30hhU974/76yLzdqOTF+02nI8Kx0q5MYD4thkQ0Hs8BdjC3nXLgrSw93pzf
lZEQSe28TYSrie8gEsUJjoeTr/J5W3JW7bREXnbm3q8CHhXZW0KuLz8xihvh6q+CAaqqk1zCi6In
Sgg1g4FhqeXa4VUfOD9KOOqf8pSxE16uCdmAOGipbogwzf1Telyv3+B4RxWSHqvwbv7p+j2yf+Kr
nC/hKJDm+RxZua7xs7PCFHm7eQUG8Xur8rj+3lP50hKDN6gt0SUK4P7B/WNBDvFLTRQgoQ7bpc8q
bobhranpWWmM8atQ6GnoShIPbqfOgAkJ9gItdVMSN2DGpDv5qC/Oomjh07TMWp19upFMRMi3+6mq
RYkzR1r00Bnl6AZpN1ax2NB+Gp0De9n6hGy9x6afqci8jOxtGQ/GeyfYxQWQlQEsFdiJUWDDa+lB
pBeDE4EGNZP8vKeNMZcg810tnxuW4BAw/IOGLBPUXw+Tcvltiy38A8+2wv5RMJm3CiB0gcWPl8MY
8QhxNq7bwlPsn5TaBD2wRII51oelpSGlMAsYugKL+73Ovdbeb9txJWzT2I25YWueNRDp03eQ2Lnk
JETBc5Lsw12L4wzsyvrufb5wfoDIgl0WU+81MvMxp9v/0TZmIzggl0tjC52ofZhVa40kheNYDgRQ
h5RProtJ/xvq1b2Kea85GvOCymxwFaRzSnI4YeMReXzou/g5pg4BK54gNGcXIXItZtJps7yR1dj3
s51hvNez/mpxFxb6KSS3zIIVfjfOhcHEG2RSMzpDg9MX81KFOWVBegviKHnrj1BsBE8S3kbnD5Zd
3/A+Bcy577RYmOtRj1vaj/kXGXv1gDYx6ODlMeUe0Xhjae+RRGvqWzJC6V9coTGCyauJp0RHesSh
1MYGBtdfHVorYsFt/+bmrMcr3zIPCjmfF9z6oiVdkrziAmfgg5YMPH8/lGCu20GUYSrJ6axTXjJg
J/bPCipWQh4GDsypgOx090CfUq1hhNTwgb6hXsI0VGoQvAeASYCLiE6s6dj9tcQVdsmTcPlOM2uM
lRY7Apxi2UJrmAQEJ3f/HHKg+NqCuMobt42FeKZlqyL6wKm2FSJ3zRBS9VP6MMqUbSO4p/hhhE5I
mG6hrGTd/Rrjki+UMATT2XVTTll7kWy3CGI5K6nvdBmm5WbDhF37ULr00POZJxr/GxwOCsqNm3a+
FxoVvO0joW8IrZs8akvdtH2cY+Ze6vOaDUC/kkDNQ/RLll0PYckHOflPUSl4T+6RfPXpKl2s/E+V
sgREhy3hhBk/uCBASt4JesDZcMrzsd/gfgF3up/7jg1kaOhCMAtn1eOZq7lgdWWzNpWPxzUZe5S7
MINK9GsiysI1Ylo+VUQby03x+VM/OCPHhGR2ZnJkwXMiKuoNHL+RrstR0d+A1nU585JZMSo7vyWE
2X0iY8MwTf6pUEB9hr6Obh8nUqBH+7stg+ikNm9AOiazTBU1uVE0MsLN+y6aBEqx/qbvtp9NFUqZ
Cpl2GciQARXhUcwn5xn5ItD3NFE4AYjWi4Fz/tyEqJI47jqutWB1LOq6ubLMrBfRADa0hRuF22Zm
hTUHtWjGbDgSUWdCcgV4jdUtf28uxkPbFyuHNXRhsXwAW9Tcfw+Z9PeYec5quuHx3xjbWLQJZmKu
kn5hcFSaLBVOU9Z+IWDe/3pbTFWP2yevwP8SWgCWP7x9iyg9uw9gbfRcLwx3Qk4d5iaNKUS/G6cn
D08oJdZCDWY0Z2ti45Bpaqgjpz8zYTD723MMvokqO9rsjff+gtZ3JYYpc3LZTAN3zBuI82/x1V5K
xHBTU8nGvxJWYy5O1iuRPAAkr9HvQnmlFhjEslZkvytS417NjeyFEuqukVve6Na8ELBno96rda8m
Ew4K0laE07ptMmOJOzWr2SIoGWF9Cwf0e2KTNVxQPRsO84ucHPDiUkDGo2IlyuWTm7R7IcKqPceh
6J1lQEE4JCebpVqUuzxAhcWeE/HyClEaoyaaB2I8EkpeISzTJKrnsmpQ+4DoqJfAYPLU11uhH0gv
1zb3R4nynNaSYNyV7XSWx0DigjgiJsluZ0xEpkGmFzcf1+uYpI5R2vknCAn5w4GSGncx6zXfyow9
SwnHRmuja8nap/8HFDEU6zxs7/47JPmAKtrQbyqYaHnrwEyo+gzXq3Zi+alQe8ZIxM6EQVm62O+O
W7HqikBubM+1BkmvOlXhVpm08atXndcWgmX/8AtAyBVALn2fJgUNy9cPryA7cpVDfb5O+sjxs0ke
A5hZwHsWfWn09Dft76W6hyrJXYGxqkH2JTelOwYve8s4nG6pCNQznU1WoFvao37iiBriCs92oxQY
sxe3B3TtnXokOJ2EFSAr+28Gn6vJbCEZPY8iOYounRd/ZmSN9thp4cUyC9IsvHvjQO6W4tD/qkbA
ZliIAMqBzAjdm9BnCigxeUweawBtLzF9uLQeUknRs5J77k8RkpXCTJFfbjTUinOms1jh2DlmbMxx
nnaGlbetGJqTwsw6M5mCpujwdsSRYNcIYL4amxvRavijbj1dSg5SRTNV3IUEUvxvpe4yv2IZv+uL
leDZeubMSJOVK6IXSuZDI1+Jk7zjOUfj2Tr+/YTPTA1EUedpQrcMN4Ynf3hzC9kYHFRgxmSKHqg4
Gd7XzIf1weFNhYC9iAYf1aI/GxrrE5W363XV2TDnuUbJJ2y8jISFV6ezSgCatb6+FY+5UBVchTFi
d3ET1+LwYCdgAX319BmHEJV9blcZgc7dIBi8h4spkn/XEu+qoCqjtBTL6Cfqk279qtHQguhz9Kkt
KA84XhAQt0NCns0LLl8m1M5QdibjI8lbiPaI9u6duMwE3trg3qkxarhhTrdRQeQkpWI778Wn2xAA
oxEnCiLMlG00tj3FgTvrlY4n4qActIy67e/tKBncsdMJ20sMrA8sdMwbSFrtI/bUAESbv/Gdpmz0
0meaF4SFF216sd7ojXMGl2vCLsLKdRrZWs0Ykdx+52yB7SaR4SptO3k8AOybJq8ANMcAaUSYVQwX
BSCLCsf7jKqjVmszXylWGzS9wRIGIpJdhfYWpkGrU15Qep31GjLClCdrmPaSEuVhRaaqA85hcJ/g
Eko2cct7tB3YrnZ1oSxkwNIZB0V8XW1flIaTxiHuLODvccVWW8IwfLlpBkRTXBBh/zCJip0fgBJs
DpFfFaEuuf/wQy2kcXdx5PvH+gXJDbGFCtYe0CpYYtz/wCf+o2oE/389DNNi1hShdh/UNXS+zc+4
W0BA/wwem7DGReFo0p/QpoNPgCrXMBIoYmm9z9OWSV4uG4T8AzlnQe3EQAgV99WvYdBwj1hOW3aV
aNaG8/LpHZSlTSUrsPSFYeDG1ghUFBSOqz5HTQl+bFVyuA92A+xGB8HVrL/C917GpAlgSevS31eZ
wZkFu608tUN1FAdsXmRn94EkkvQAW2Ybd0iw4VkXn/UEjUBdQDUNwmFNTedXWYdtD5Vc4Sflzqvp
mV00t6ZWi9BJPDeqgzHh1dP7DjnvlrEUrE/HGdMfrlgzXLenXKNP7EFtCJB9uf83/97URGkUg8AB
LehkpCSC+pfZ5oBHyC1suH8cllcylEzrCQR06GUJeSH0UmcgT7uyrZbhIb8j0QW1J9Yl8YWlk8Re
xcVIp449EFTBaauoRv2FJt4fMKV9r/Ujl0fZjO56PAgdEKZHqNuNatrW/3gD9xGDgVszojkW/B07
y+2ZH5/ysRTKpfxHq5zGOZv6fXqpiphzCwRqXh4GElgNmB/9+39B1T0GTta+/ZacSjk2g64qUlNm
QeZQDxK610TljS8Oith3Lc6VXCkr1kY5LjODirA3MPOpzkUalQGEHk3vDHKPeZSdZOHiS0Bmw4iQ
ZXbsrXtK+UqryFOTaCE8hHz6WP4KGDzptkl7cGYyNeIzn5BJ7+2V5TKSibqAaMqU8xnHXkiM+mLF
0YyI4RNTvO4iiN76uldVQ0/d8j9VujgGZ+tkEB5R3IW1JP6GbiYP7iqhIp/kMv+IxfhhWQEe+AFw
3oj0prl59NHPSKRqJWYs6+JCz6lsmXTHrhc+bwNSI5Rg9GH9FCPrFB0KKwWMtblXkAbnwP9+IYFB
FGvaiyUdzZdtyz5G8HPFPl1uDqOr/gCXpJlMrgr1Mqnvy+4Kasip+NaEAWDzNiRRtT60ZZuyR28d
DKCZE+/eX7ngBeCigcyATO7sBnc1483GUFAxX0Trf6cMLoSaecL31lrXW7PaxIO0xF7/3d+SIh01
yIZX/7rNfDvbad8wgzxFKQtn85j+t6GywExKrq/dLAz9rTMBI+4C5XvChGktKmOe4gyZo0PZMtfB
8fCebqK8Yu3+7a7puoO/jl55altdTFTATYW3fdoobxt0XMmNSukHduOkfzKSKLt2y7fRwiSTMtVX
NchLgqC8hoLuSANyOb+bmx0UuZC+KCo1gw6JZUbwd/bMpQ9iksGiv3vXBFw8XcnmVnDYOPoFNS7x
CE714d25/f6woIl7HM3EsyxUMO+3Dvn/c/4QQMisRRa9wbUuAj4ykYH+FI2E4h3hyaNzp9jaFfuV
wffayQbCyMxDDUAWx0uS8hyLxL4ZXB6MVnjDO+1a+RXTFS5zO9yNN6mRBZHHN7XOiFWgYPtMrhWA
oFywOd/6qvNEaTWIgYzkdhVQGZ9gR7UBrrA5xDdfadKyFAn79t0bij4DmFbQU4gaiLU/qAUQknCs
IcIKzMv4LU1eQtzf3pZ8SGWmUfE8VpTfGrV8M+eSaQaz6E2/o8dPapw2zjFAQ72CnCD6C5B6fXBd
DW6d+PAirG2ogvQF/t06VGbFBvpgTjdnTqu78RXf5eV9zc+vAJyZo9mKxMCIYHKaw3Ikuo1tHvyq
D8+j+rgQcXYCTAGpajjQbL45zxVoNReTQ08dRRojU89+s3juS/szZQ/G0gSCw/yY9IzltQPXyvaG
3xHrQypVLDwx/zzKhekrMRUiO7lWqojRzsKNCGfwihW9+jfBPjn+qYURmM0lB/waIkKWAHMa7hQ6
TrVJjO7YJLT3ZqeAYj1zhKFqPbk0gnGF1NSYWqOFsAeUGjb5iXPFRmB9EnnSZ/hlNKd+kndOlBIr
Ljj0mFFEXP5dYUMd7b3kiegFb5yt8CXPMkkQLr5Cb8kpT4/tpuBuXJQAhPNUlT4aoi7gyRwBm8W9
p4SPi+a8YDRIGIQz3NAkW6+nJmzzOGFHXhUEEnKhB8dLlntAqDDByllF3nZaJPvMxSFd2U0afEOO
GYH92eQIWF/b0hW5bPLl9snAnfF6l3m56nMjof9/5B20uSfdVFkj4Dxzyq6bWTZ19j/7Qln/9nRW
ymk0tGSQGNUHo059KXDRYs1WoK292Vcmhwqn8PLffpURNhcBHKYX1nQtHCzFiRz19L6JWxro6Xba
Ucy7DH7nmvohESs0+w5G5rIMOSxx37T8kYV1wFF4No3HAQBszc7of4VkmC//U+q5dlsb1D+GHbOI
/DUPNSAIxMs2MONsoTnI1dLsiSd/ngsqwiS/xD6R+qL4fWI1tw/CQftth/O6Je4wsrU6qd0v/n4+
/PPCpwNZUg+Aj3ZMygj0SVhvxV7e3NV+GRQw//MSzEeFG7EAhUmo/X6Brvhe/TmNJaEqQpEY5wN9
XLC7Gq0sKe0UXscs2Pzk2ULIrZqlXDRYqpdaT5hH2pix4qAmvCw+xELt60IU3z33RGqJzpdn8xsR
KJUwMECMXh6jyFekXEjC2G5Rz6hcrpnapVreRA3lJJIzobqWv98U0BkEIIintwcdRsUH3GOhnptG
ycB3iyx937b4IFzLpnDEaCkXeKCQvIWmWUFtfRDq/9UaGqvp6KKFZsgRqxNrYk0WCdbKoVxRnA+L
KdHorzGooQrFLZrhAa7mKmNDPXZyPlSeLZJLLYDGXcp1MlMMimNzfc9b0BOkOaGhmPGeQ6CPupFw
rsm0N/0E4E5nC9cNnMtD/X5dwbwGAbepZ+SYChSRjYcpJ8P4OAbvjEMiDCOvb8nwyYZDPE9y7rl5
OcIyf45yefZsVZvtS61iwRab7jpSJdXYoANgoEKdc0Mka1OixFmE+eM1Kon+VuaN7w03iKxxHyIa
Om9vZAmNkw31q2ahS8r+e6uWJcN3AGDROBCiG8z9Xw6siRWxkzz6kAJ+FFLg8f44GehBisHLFLT7
Ocsveg8HnoF9Rvm3ixzvBN2Ino3XC5iJZrCtKvImQStzcuQgzASpRLjm89U17Q6H51s+i2fwjjNA
SpIbaPoG6zTfFNUvSqFTTqtP4oPQVtjzkpbzFYOR07D6eg1fsEraOJ/9DIFtTCgzVbKtXVFa/bhv
Ch8X7ZThRdQoWajz0FOCBS3l8DGROGDeHE4j8TGhzqI8yblfrtpzu//7TLmVJ3X8H9Bee5gmWpCC
J2SeeQLxGBEI/3+WbQKMnsPDHmNSu74j/4h4I3TdmSVqJJvu25kOdEDUG/79t524q+WoySnkR/3K
HLLNehbqnKyd5J854dLNpA0z0iMXugzUeuOUqEuIvSvh69HQgUkvJhPtEO1/PTB1Yzg0PGyZrV/z
d6pG3Uq14v3RCR0d+JfmGT2PS3+OWeKzX+rAUan0ycM7/30DSrb5MEv+mWCMRKtwdacur0gmi1zN
dtiXGNezBpqmVHmnaCxnrfirv0cJhiUJBWNgKNED4SgDwSG9o8y3ku8BsUZNd6+dg1QOqekytpRO
ifDVYH8PNHKlD8G0zn3Gd/VlTgia+KzI5V1QvceR095uJQHfytydqGz1T/GNe/QWi0rwafbB2VPw
7VHq9KhYkVUIGjsERYFmIes9+0Jjdmnz2wbjYtlqzkOJac30h71RnhtOQt1Rai0YNoBSmX+ith7f
5gDFfGeLGt7HcJ2JUrOPSpTn3jScU2dZPKaj3uLOdKN9PANHfsyy8ZN1uQL1pfcAAAJ4AEhr+Fzu
pYBT+9Qq2JWrEHVLi78TjLqOBYQcjUN/0Wq+zGQd3XofoZi69P49ev9AQndj1tLKATw3T1DTT9Vv
K7dua1s2a5XYGa55jAGkkmR1+6kHg4BzOfeaaY3Mk76HwskVd2hHwSTHAclDxBh4pbJ2mAEtYtF7
otviIN1kvW86qIg45cyaQto3p79qyUtM0zPcUEnuU5v+72/+pfyxpwrBbYWIoc8ApKnhpq6Hm/Nw
Zbe9NEC8lQUm01YPGeVFM57zr24o6ZCd+DmzHx2h9LE9/zznsGXgs9+hySO8rO6iwR4i/dpJx887
aXVMwNw6cDD4PhFLsSUWmyyrzX2+VPRiXTRb7zDVjehMUPe4aT1LRpX3yGO8MNDg0HXGk3Jmd6ii
v4KOz8s3bQ7svL1MIdxD1FWUYSlldRKei8To9/QuixJuRAY0C7RNOdIKnEdETaMqL56mLNRpLwlV
dWFIV7EvzsHfG3CeT/toYVOOEez+rWuBJWpVWAYm+JySXjq8VWpjedrZZvofYBL/e+qxQmPsLItC
iqYrGicYpHBseQVsNea03AUJOtQvRwsI/stjN0qrYQ2Ha8DdK+ppmIn5LBvlzi0L1nxYzSLOmYRC
XfYkY3EXJPHQOITFCpB70pb0YiAgKiFqHs+likOYh9UuYFFWjzsfraXm5PwUkKB3HrqXKjFwky9p
ghIgtJBuos6AK0Nx1JKNnQCgVA5XqxEstoOzpzm5M6XY8Z1iyH2nEA0YN8pcXgrXhGf9sl6SCpao
1bcZj4hTTrK7C8+DcRoMJKMOeTvze+BByBUwdKL0OVEFIvMwGxScX6KurJvuL7Is4vZALPhhCXcW
kA2hEHFVhCys7vh5IVFzlbDeWNPIbCoAh4D61GgduYlIxIPhZVtr+OUzySgdX9Rlz0GZEpSxFLSc
jJjHuNJInX4XlyF6JBWUcz0NXJEUMsfq5B+k2paKkwxqtvWWEtu2LTXPILFFHFaI3sAABevVfp6P
ghfGghvOokLsYXxoDY/XMun1+pW8ItGuGtijLOyTVwVp7C/has5ULIFl7CqUGZM7uebmYiD/5Df4
onM6BXpLLPAhb8iV/FuB7Hw6c3s9YmY9JHKw5h3cFXNRTpBFt0NKxwqdcJJ8UvroDPPMtzg+Sem+
q5wNBGTUOp42+ep2HU5iVpeuTKw8SLuWEvUCpXup8nVGrI01mbLkO499qR1uyD+BYQmXKbEWPE3S
2Ul7E8NhHlsGd5nybdiTtlb+YwX+H6td0P2gh9z67Xh8Axev2D/XZJnwhNC2Mj4OcDauUo5oD3qn
SGe1k0l/Pe9fAbN5d9XEVH1wagn7+LPFfZ14aV3iKrAtL/kkYTHxh9zmPoIna33R9Q9t+Ojg/VXk
XKnKyByFkgcGmALBIyAHYcaysOGuCfhU+sD8iWE1/NsTGTmLzJJKQT9s7efoMv2+MNmr8Hz7vViV
i8ot4tnyJA1x3BVLFdqal0boApTMgF/fjc1UE2hLn3kFgC8+lKDSogSsf+IKjTOnqrrrSOzEirfy
9q/O2uCxWb4vRoeoDlvEH7qRh+PLUlfCouMaYTdvgvSjOBubWDh9o83ye/chrOL1TWscEPhjBatq
+2uyJ0v4jGY+WOSson3hGxHMkk7w8/PqBVwAVuXad4J9wqxOtdBMQRBUjqdTxYE85WDupyIA2y0v
E7UF46geiaZ/+PbS2lpDCN7keMudZzVNY6ZO+0GJfrGjGCM0f/J5GihFtYdDVXXy1N+K6b80KfrD
3sl4VTvToL9IYGQr7EmpUNx6ZvjXjvLPIkqv9RozsxbJyYV85slU8ezk8LkLGDZ4+QZsdptwcRJ4
CbuurRbIIFRGFcE5IjddWpNDkZ8RrJ/zjPlm8rRIax8+HZ2ukp+H4rpqsBF4k4buYly1J17hj9sX
WlEnXkxEQUg6lFRBygFSuyTSELDIEgwre4n3kqEx/tUvxbV/Kfm9To8/6//GKVyoJ6CCR2M1Wqv7
QpR7enUphq92Ordk9S8ABngtQUhFRorUhTMPbb3RgGAH8/mgoxbV+sX3jMZyi81T5tUleLruXEAf
7VYBSSIHtMAcGqhAngJu+QrH5HHlcsNY7+eB/+JeolZNjUzO6xx4obt7PpY+HMiL57xkmsvjmwTf
rWjBmgPcmbYVqdeY+7DNm3Cx78jf6aHyWm3WsmaQMHCrhc5QbUPiTHEv9aE14+IPxuiepp+VB2mx
dJ4nvVcE19YS5gz526kfrwbiU6jEX1qxtfdaEjEMkHS8ldd5Xsg9TNYYnQW+cokLd3RBy02PgU4m
MYIc0iF4jvqM9XKdjPimGhASeZY6I1Aw1L0dK4TGC5hRGQhzj/xn/MFX6bsvrOreJgj5blsg8lqP
8ETRrYoE220oGUqCqF8DwjZHpk03AdzuKHtlEpCLLMAeK1FOoj1vep4Qq2mx9Auq2cxp3zwlKQa9
u7e6OfiRj06rTjGiqUfdMmHOCL8xLSIQ3FPeK/cpDtNi4iMdYIdpR/IPNY74DSqx0KDYdGoOdBVO
iSUqSzIexDVFk/yyBKCzvvtERp4nHrpuPSwHMvO4IVaAnoSyfZLFJ2FcS1difS+reERps6RaNr8y
b0htkgmzKDczpHIwTolJMVk2webzCoy/sHIeiIHSHFe2NeyUTo31sYrecy9ZV04XhdoyrgiKmkqJ
Qje6fVdgC+t7gw1n4rGJ5jvG8r+5FX383Xdj0zcgpYIPZn2ylHvPCiDzuPmIcOAYjLy+ww//i3NZ
Bh9dw5bg6CYsDkLmni2A8+QPfAXZmPhCD4IRx3abxCfWaK6z90Sm4Fw82gRvhNwYeqrrihYBAkUV
F8Vdb3DExP9ZKg1XmaT9hwA6ioVCCAvWn8fSA4ZHaiKRjEa+iFe5IJxIig3hiCdtmqJ+ufwaKYtB
KHPiWY6PUI9lbuwp7UEWSy3xWbr256JDIl65HgAx9Nq8DSmc4NT2GJUkV2yqGPkEF6qROqnLUMUt
7xwg/3/9yAO8E3fK4+k1KjJo7/EfO+n8bjS7PqIXa/E+YI6J5PaNiHb7Pm+nQcKaKCq+3jdXODXj
kNCQqvLC2m6242b/O+pbqX47WH1VWA8Sh8zFTuRfl8e/7SJl7d3/a0h7vB2NbFnxYMwidCkEx+C5
XXoRkRjPTP/nuvvKdtF0uKOhE3F6sLo7E1y+Nwtn533fsYL50+PgFSOsu/+D0bt2GdIE4GVlomNp
Uk1JmppnsGg27RlmNdLWtcCcdSMNbWobAdcRmkuEd/CKzHycdRHZCbK5Yhwu0kX1pzxNHyDL0cLB
NV4fuVS78BkLe2NSYAzHk5+Q4z8BMi0+tT/H7LTVAavnUBlDnN0AdqN0NEHBk6m1PGTD9r9s+Pc5
8T0JLYvM+hs/scY/P9j8FdxKukcmLzjWlBZTPbXZWp/Jq0EYmS3Z3aFtGa/H8rRn3VEOhYBK5ofy
4s0R/kr74DssDA2Bw9F8n5WJdxrxS29hj2gkne3GCQZJUXUyQ2Bl9ETK8bmHMRdf3sRS0GJrE80V
SRdq38Mg+hRTds8W/q4Si97l9fleo9mGNXhsUsfoHfJDhkggK4vXfZ2o2h+Qm0TUW9q1vuiJN+Un
qqBm/U8AiYEI7pZ/o5oT80f+R3GgjjsWNs0Q75LPcwFl+dGTDzJPLpBGV9aI+mqHMZ5OIZ1uuMO5
QW83ipC+Hs+uC+gXl7OBmbX/53MFFYm6bfRYmcPgkdDpJXL+WapBqoNiaRXgX5A4vnim5U12R02P
sQh8SGlIfJdYb3paBYTFVi2vqvhJWe62MZllnoMwVyF2Oetm+UsrTRgcTMgUm36Fwf02zcISicaP
u/ydoFNeJ4DFJEXm6p+J9fY1J/T8HFM0fFwsU6feA4GgG8zfcK2Mi58A/SgGISr4JzKmI3LTJQ5m
BgrmXO7wtr8BnEt1h+Syk+e7Q2hSCtOrIHyljhnXdUye3VbPQdDdSFfWBVTxNleASHMKk0QRLXFg
olVhFLDqdW/8YpanwP9/RsMamtBaBm9KKFzjJJCh9PpKS6kp1lNcEBpZrPPLZ7L3VTVGYTP39HZ8
PtHRNpBC537nvIfxcvvlBcgGDmEn9H0MMMw2QKCnOInqvst92lLQ0yNCOF8okz3zVilcZYZNEGYJ
dabSo/7+ak8etCH7dmWqni6Kyz8IIZX5k2ts2rxCm4kk7RvU6roJHu8BZ5mqjCBD74T7gc+BtvKf
IG+B5Yq0sLyVS9yknNkSLM7gWLJTpJzjvuEGqG8rNY2y/ZAAYtadDcbFJv/mXNoZvg2d2bGq96q1
W6nM7iAmANWWzVVLynPkz7PEJChiLIk8TLl1GMELVhUDemMH+3zjhDQRaseAyIXUJD8Mczu1xrPg
cLUH3TkqNFhrczU/C+d0rbrw4AkWk2n2PYrlkFAzTLduPfSLMwXQhkhsfvKGvYUAUuHIGllWeq1d
CivCtHnQXpXQqA1mRtJdcvtY1o8aETu+ewYigh0BULocqKX8cpuy9+nqSsI+PaIKdWz33CsnIm1C
icp24ChwicfRkMykT82y5OL2QB36zsFb+TCmZ7f4YsjTeGwCZleFdvDLHMmVsErcemhjp+xifmJP
Io5toCmKA7Gu0RKjPRkNiMgncINO+A0xla2OubfIpRtRsxgE8NWZ3w4o1dS4u4cA8vPC6YQuOYu1
tZ8THVoqHkgUu8GMjTT3gXScMCPfbUhNYwoT/BWNLM6aRjpoqDPxMeK+lN/p2Onpg1V4spM/xWwN
jROCdjLtWee4SiP0sfJSqxCYI8WUyrp/skGtS+hEX2Ag5BCjV8G85GOOJmxyYcGohj9kN8sC9tOL
DPVxDsb2MUpi6Wsk5rGPVbZx/bdKZVoGCqCZEapV5/VBSpTihcHJ8fchgL7gHpK/lEvMJN6Btp7J
cHNBgCTCiaGrJWTaUOk6rSogDgWr+FFxpaJp6wACU3sm4EdLmsyHWwEOTerHfrjTZ4GQ67Y80Z2B
qGkG9ynQbEla8XzHm2We9RzArzx/SWcfnEcu15qvW1Eed4Gs1eVbMwmRqxwme+WLEuQenR5+u+Hb
JyMo147/8aT+oB3pfw+verqpOroSlHSzJByvPJjK0tiCNv35tTS9Wa9C9P/g4eWVIAMeO1jqzHiq
V6WwYlnjr2pzAPKuVVC6j9oe69aShgFqVPYNVEdqNLRUQRUmRhtXCovrFexWgE1HXkKjHjChcZB1
mmsznPsE6GiVc3/9spR3RKFO8xLzx+7ZJyGoYbL+GthWPMqI+g+RjWq2SrakLotL+Q5MAjqppC5y
Ctl19xM++LywblxUfIhPlmpDa3EZoakpA3/A2UW7V8FyHsqy8Jmjs3dp1H630+AralC+4cgdbQUa
ThPFPW9qrF910LpRS5ufwwJ2qCq1E0ib1bA7o6lHyxhQSzFT2GYQH7b5okjt8E39ctUfI89yVlEB
r8n+fB7Hwu/Zt4Zf7Quo8pbWChZytRvPH0G5vsDQwCex1mGlQRQLnVTBGt5+p8OUR1hTPDxdWAJM
Hz8VlVFIfGEvmVN2RLV7zrsyTogn7JzSD6TAvTdO/NwwmKzGSDJDQi92nhGqgWgnD0rlSRV9l4Fx
cD/6m1Azp3xdUU65HB6/Ulk9J73GRj6syR96sTEV3qFEj2BzG9oI4bP3NZiuC1uN+29IwwkzTilF
ln+eoYwPVQg0M3tcwR8sGduaJhFFOxggiaoVagEmNbdQ+OvGY6Ob64BOGf5N+a+0VongbteoP/dg
Q/g1ofltzLJW/wIUp2eGsaq4x7twhtSQm3mBileRYQ9FUmd4P4hIcjHl8xxp9kqURmNHzqLzWIwu
pxfEkiEydk69q2kkjPy7EKCxP39RKjZsuwgDTSpDF9xWD1ITs4tgOhK7RrCTTqFmq7eI1Wt0IfjI
lA1xZix7LLUlDDRWIEDCHHOTWnwhissXCLYeKX+L/XEMNeob8pmeoPPnaunZjUH+aW+89AqpqA9n
4h1nX+MxjXtbNElNzEnmMYuROP5KzJODynfZvpmE5PgVcBb/02HliOx/HEEWS91MmscWDJes70As
VR2m6loujowdap3CIlAqRNVAhoQ76MNrHDdgjaMA54qVlhZGVcmS/Sey94RC7x7LpGQ8WG916+uR
LHrxJ6uEO2AuM33LBx+h48yd96mJnqJXQA93qKDBNNDjw195pTI5TGrl57jhur2muebayItADJO2
qE4m7fwT0aJESNzUHg2BE9yvA24Jt5G2rRi+dulW5QmvcN998YndA8GBsWjY1jY9aTCP34abgede
qJPuhHdgwpG89O2kBjC3/myresONonA1ro2tthHjTK5BcKD4+srDDczMh1/wOaw6xbAGSojnkSjT
WQ/E/ywSSXNstXtujY0Z/h1DaNcd9NZh2sUrq+OcbJ/gDpts4i9XSk0rgJewf1VimrA8px2TJRWx
6dZ/c97fD969nndvDSE1tDY4IGucUlu/60nXyf3SJRU6u//GLFh9jFbmvJKHYLVyRqJ7SQaZttSx
GmTlAa92MRV9+jBlNSURtJTU6zBqR3UVOoRIgU8ZJOjcFV1XWmR4g+MHF4GoebGQF6R8nhk+dDOG
pi5AdOaCJUQO5XIaLj1ItWIAjY0GXdr9QFd3y6w/cLKUZ21wtzTyOP2IT0WYyI4cIk4QXyxkFdhi
rYtNRA8CbYH5eRcnnErSVT9b5xc7kjdHK0t3Goqr0DGuBE/8jIYFnULFsRazbTpOBDFc90z8F7Vu
Qcyb+Jyb3FXZ3hUTGpO3KI9p/QYdzJI1dkywJGPrlDY2d3VKDgdkJKH0drToaaiDqDzAR+CTalHA
X0p/3Dyr7/dPsVuGY0b9Y6CqP2SUxZGVzRi4ziTBtKlggPRNhwOcOLgdX01LwGirjGDsdN5r3w7C
/Rg71HO0yQel8mHmFgFgb7Hq8/rO7Zqviu4sTzqYOFKsBSNCudZzVvYa1zFuSqiG/oktLiURfE66
64I7Z1U7oT01wx0F/0W8h/UmrhHG4kZnRu86Ds7xrhZd0mubT5lR1ycAVt2zMJ9EHjn47hLtioib
XBjEi3JLapavxbLsuVJO3Sm4Np0rvdAHjTawsrutxcVxSABL/1GEvPtssoGuE5p681yem5ivK47G
ZPYlNQZbi/DWJ+UfTWQvi8x1O/J9ifMLsS0osAzaPeP64xJYtrz56qKSBUGWesUyGxAiD+avs6z/
JSwY/guDwSntvXTaW2nqdIPNHlURa/AxTDNJ2/EI9NX+/M1XYaM6s8ubxIA2J8aqjS+I9FePJCE3
YxINxb8A1Ogdn5WObuvnkD5YMOrvpqjzb6PBnqZiLB4R+sj8VvLbJxvxJTCvgSCxvnaXiAxmv2J1
mFi3A5wFCfruY744DDtaLBvyVJXR82QA8PDbNTQQbsHL5aBIIrksaiXBXZX19Pu8z1o2udIiTHoY
6KJ58UwDGF8HHSNVZCWwt4XHnc+bFLyncp28v9gqDnB57AHb6uwEY8xVZ1kTfSLMbZm4lKFY1IJb
WkWkRK+DK2SEI9qjmCANXu81NzEUJTymM8CIYJF2Sw20qNLh4henS3diQRuMVrXBDYph04LbE7om
NCqKDgw2+RySBvxUN0bZFo5U6sIN836/zmKG43mwW0e0iHcAgZyRFcHMo5ccHc0iqZCAjU//e/vK
Va/lPazU/0OAvxhygjKwhJ567UPvQPfJyV/2VopaMmYqHFqNGbrV3AQih2HwgZ6pdZ/b5ywCbtvD
OZXzaQKnK0nXesGS8T0MYk4BbKHyBrC2DobdjC662ZILj3VExlqnjSZxogRQ26oR8/ATNMcUUWp9
UeQmpvgAA05GpMlcfMxCrRWbf2XObdhlq/NSfIFRG5GzTMzsuhwt2+Gythk0WVzZGEODrrqgyuJ+
mS/EvhqUANH6MLNfWxjSnrBLVBE+Hsjt+zzVnXGZWwydmAqVSqPdq6qnO2v+5PsD1LA3wuYOgDID
3vWrfk43KtTiCwzQ+8wGUkUavFx1FFnAH6zsL8KTLB9Dum12nY5xJWIZ8tniJZgRyB3B90H1m/XW
njB8G54vgJPTe3ivcMKFvQyjH+eSHJcAdymh0Swyriaq4jQu1JtA19ZC8UtGvoc7Ex7tq9/rT4pM
XWKSR+tDRfonvaJEshrh67n25Ac2MRy9nOM1doUDl1YE2iJY+7kDf+6/EvzMxBsDNO9lcOGACcFF
/+3+/VjUErCw1T/KUfRsKG2NBFQJNXNs4ps+zFe6ZHyue5cLgq768ZIe4C/mYnDj+BJF2faeED/a
zjuGMr21ATLiAUv7DP+fHW59fzaKz50XnkCp4aukYe6tzfMEFmn079CMBA8ahPT0r8H0B92aN+cK
EtxmwN6RjEVaj4eEYlgl2Hsa0hlLnd6s/QUP8OcdGiHy20DICTdqrESQ07KxFbyClBzWYOK1TYmW
TN/oKemdePhVXCu+v8edkrxQ7E/8h1hURt298ItX7q/Org5aaMz4BsmzYQhvVBXNZhzgV80n32nz
htdBm4Op1vS+EZjBm+Snulf21yQtilyeGKAHCxmt7ROi+MGROqlAhJDFYg3NQk4YHfHukseb6dqK
c+eS0VUwKt6Q3DmiPMg4W6KiN+BAU1QrQlipLz3XEI+3qt3hTqrSQLI5UDy3jF8jM/OGbm9X/3Yj
RVl3mB8tJtoTiipgmwyUnW8YJChSeGhwGQ1c4b+DXxGVjrmlV8DG1M8Fe/X7vO3oS2ZqgkzB+idb
/qc9glSbgSZgLmYMoQsRjFX6ggWRz3qH73cbvMNuMHfYjo4zmY1p016OWnt/cH7D7BFP7nWKiF9U
nimlcY9WxhsQ2LPVlO/x5w1kvOzn5xEVJBhkG/Tlx3gjv/MfNRdwlOTzfRsC33Ts6KcJ3SQmbaTR
ghwCqmwL4cyZ7gERUeDHIVYlYPc/oXOHzpHogxU8XPi+WkOwtlauz2fjVWiR9jISJs9tuB5hGyKU
RyWGkFMMUR6oKubgkrL7OOIKEbUxhUVXLNwlUyqMCbeASbb6XZfGIvp+fl7BLYQOzVSAwfpc0XHw
wcFgrZAL3NhNnOAqV76LUOmmv2pYb/kJcSQVjVxvZOD7O6RbTUDUnKXoVlkcxQvr6dEwSlvNjcJU
07+VpP/r/zRGpTd4hpOdvD0K9ErGBtBLqPQUQfG9GXiUd+2zQizJSw8vFtzzR0kWbzhuB94yPE99
+kn9JKYxlOsrvl8ir4ylB8WyQqjcTKv9p3Cf1fcm22XAR4ShZmD2rqwgXlankqipYSShIBQyHChg
HVFCoTVnVAt59o9CKA2J08mOnZ96QSIcLBwWcSirBZ35rS0UzQeF/u5poyhw8ziSinJaojxJp721
mIkcZTiIx7kNeP74/3SRiGTsaGwf6Ni5NIAl9dV9PZuKvDj9kgiFPhHmDRSv6DSNUnyEk6txsgO2
ffoOnbL6zjbcR8RiWdBM806LlURcu7mwVpDd5VfqsRCgNSc34CcVDzKIXCppXN9ECh7RwWHY0kIV
dq0DFxRXZLV30xJH5OmlM8HTAJA3EcX1g7IO1mQzCQrJif41b/Lvxx8/Dv0dVuLtkr0swOv2RIA1
cHjvQcOihyCAgxrSmZuzC7NU8W1SejDjEAtrj2ByHo1n+KCYfebgFRyGPXS+RHLo6cPs5ku5vTdk
F6LG8dpsmz90sBnZ7Krw16+lh0FfqJuaXY17U4dKLVKpl0Ytu4IY23TYL/EMwSX/UUYfqFiL9o6C
TwPjK4uiL22LrGsKotL6G84A39F29ywQL8md7lNU2Zu6jWpVFzC4tjZ0p+OjL5vjuA+GVJ9oiUiV
FGLHgciAWSShLNvurfvuZgnFdsvKB1GqZ1dyKE8691cbqMp/yMenlQm5AWxAWwD44G7LmHbItLOL
s9QEiT48Lvkw4DZk8rBG8/mEVBV9Qx1iuMnUT+fqX/4R7Xd+NKK24NZg/S+GjKpFQPn9utbpkmwc
ytiVHQdkS2098hSVZ8lnJn+gUgK9/cJ/LtBMNT9HNd6M5Iv9NRKFChTB2KUKzclMtci1atn/4dC+
jG4vkaEJGiSmvdkUe3nLE2Jt/KVjGjA5wB2RaTCyhAkNa8CjgJGq+h96RJAmxNGZNsVfW2rstc8h
AfO/BGuV5BSTtonr2iCefdxMDXLX4ZJSnHHD8d25fOpMUuL61oGirpRoHwlaubbuVYp58FV+qvPm
fcKp8hv+U/m+xywvh23RgebftsPjN/k6n6t5uGejieGhvXSziD2HWk08v1T9gRW/t7E8cCEBoYIe
ZBiB5lrlbZZzpCjLcSgzTXifGnOjTW3o02Z/aMT+kfFmrQhBPZoeBpqHV4G7vrXNKa2WjI+2rzrh
DJojnB0j0txUPevLwDhgH2xuf1YT3i7+i9k2N26UPbMwEV+qAAm82BpxyLyWproe5zivKR3UCRwr
YaXIGVZ0ckRPNu9q+4GxImrONYcr7Ay8B/CFBl19gznMmM2ixpJfHaJS7uyVAUG/n4kgeMmAyy8x
O+di/QUKAAoxOmCHPHzvWvHjDwbW8yd/PJQMzsPyOwQdUVzRkzJSUU0abS3U2OHs/LeQtsdvG+sB
njfoFU5FSj73bO5Jq7viBpnKT5WNmsw5b5fX2sgU8/fMBK3qBnOU14dGlp2hsOWxs9iuSXmoIJVK
TV7K9b13w/DwMalBp7iCiOsNvjH9NQNcoDY//9LUGxGEXzPk01+yCfcZOKEqX5dHfq4OTBkvSTx6
X/Q40HeNjFyxmlhSG2uoiHi7ugqyaXsBzXYQg+OHeIgD8OrScTqktNrBJ4I0EllMT1vFKi4Q/vhf
/UKyXQneCsBstkCl69+gcDV1jukEO+m2RcDChONIw5cL0YRMvR9pJp6A6l+nvgazSNFTI5M0KaSi
b0tV/RJHcES/pGyJtQ6AMPnnoCR2KxGPX2hEzitL147wTgyWKjxT10bpG4kLYFj6azd7KtDnv4Be
mcpicEy9xzk9qDBFbLspRgnO3Ybipjn5g1CoYTdxo18nnZM0cI4GLp+2F0IRV489ZfVijtecVeQv
HzELAJ+UWNMC/KcN2+oUMxBA1a4W0U7vOpiuBqLv3sv8zkFiCas/9YEGgrYFhJlPsAhdR129fG78
ItjPRnOanux8BsWsKcPqMUIXzkEcubqivGbzEiPPxX2VsoAOPo182AUgLO5sHKJ3sM6fKZLjNyvq
IRJOo+lMnJonvoLM0M5k9xP2S0ehsCY+C6CfVfHFi59W4ibtYP4n4InDMOoR1qbvzNbWJdkQhQdw
M0gxV41jM5m7Rp1ECH/bnBcWcuKwaSDJa9KqxGauKQCeyjmI//EoGUXxak/gk6NcWy9Y8w19wHec
zkPiCA2XfljEM9Jc/UT4s19IpS8v3NE7Wqmozj33T86l7JpQLyT16BsT3UH0l6mRVOaOTGf/Hoa4
//Ieno+LMCPYBxu89oyanAJzvioQfZWEVsIbS68z+rlMv5RLnZ/DW+2ojZevLSsl8ZomE2dRN0V4
DAqjsS25sA6yyqZlWYbXiKwzO6wfhOaM+tU/sWN4ZctpFdRuoima5eCT0PQ9omV6BHaMw7x4HBlb
eWu+nboXAP4UBtQyyuExgWHVD4gXzYVi5GdEmEt3NXBSiAoE44F9qZx5KU+Xeav9ly51WOt2UuO4
BNT/8IEw9R4vVggUzqixVd+iUlyc5GepuaxK/dh48EiNGZ069g5iEaN/+p7ytrGfzkR3JbDUjKFg
P9E2C6mG6H+RRjWQ+VLzR7Hkrp/zYEsJWxnpXfKjx8wFZ/TXHu0+h/QE777iBhCLMySoYmLzMEDB
oA0z8jDYsnv75ZVtGLjlQrju0HPt4RmRXHjv4aZKpsbmQj0SBrhHQlZelCy6qX60zAu08/oCfA6I
WHKpWzTojXyzdZmzJ4XUHciDktuixNdMw1Ia78xkmip9zB7lnm9UHUkI5XN0O2Y5Qh3CLMaHN++s
OYPYdxhn69r7dHuZH/AOECaroUHtb5hLIowWvj+ETfbeDlWB2vxqAw+72a0TtrP7aoQSBO8JcAK4
xVRFNKk3rbCVGaggCJr8KIwKiktJzyteUxBE7hj8zsHuf/VlcmiTvAV3wrnZ1MvqGE4IL+Gfp05J
Png0TNGdsaDP85J9lPRSMFKNquta/eHpijtNZHWO9A1KxqbEzKVT9uM+Cx1l7j3b1p+WKdAxtyXZ
xz70WZ/MOyZQnbGYTRruCgqY8QlNSKtw7xWhoqF83gvYwyDpFsbiuA/z/lwbA7Sz3iGRQ7cHioP6
5Z5wInj/E4f8C6lJqaQ7/SuyHoqAKlANNtTz2ZwDpmpQKtptacxCiGOyrXQOKyyBCbOImgTrjnT8
LKVpV/QK1ipzdFqMQpjCb/YDqF75rOKtOvLeBrqtNec3jkmUaL4nUUgvMZGnKBWcGJccfHPmsrdb
MCrw/4SO5y4WABr/d9nIw7YxY1cZfbWxsGwbBe64a0ZF1YBSQNI8g+WsoRzWLl3O8syFtfpxMJWH
u3mcpuxLIlAYV5Q5qC9PjhAZhex4UpFAhHmccjEGryYkiZhwYWg1Ag44Lv4rpyREdwqzYw2F5YYA
VwC3NbhQS6Xf7tbzv/0VAnY99oQc+2BVZF92nftcyrP6VNHDDwzdTavmvepZlr4992MLY/wpMqhS
cdt7BzExqmNWxUtLY6nlgZn+4GrRElqp34Mte6aygYdntZLztFV3xY1ruD24x0yj14nGzB6Ym9GX
HbnLGmG0EGKUweMtGqVxJ5HqHDamVdKhyy5es6YBDRwUYsz8pKKmaYdK8YjgTZBgEKkMZGXOwKlG
1gQnJe00WwmZcC1/Bk7nZaXGEXWa9nIYjXXMsvDXLbLs/8A5oeEJq3p19TftmTzQq8Q0HULC8ua3
EG30lViWEVpJHLVl8vLJSuuCQgvDLRyRXOwF3JRTbH4+Ym+bo/9bZ0YmRhNj9ObIs2SyjdNf6u0L
o7i3mFqqqf5csKfQ02tAHft/HJjXh+decRB1vniN/VDeQmdJXzOR88xGM3Iq/A3HBHl+eY00ss5F
DqyDRR7D0ZZvlbj6mbQjGJo15XHhX9eFepMdxMZ7hFHUgIj7D4k4GR1DVTOG3Y/RC4YAyswf14y9
ZhwaqAWtQH/yPCz9yUaTmzE+9BHRgSaqlXRlJYqSffHIjRhUD5KHbUsR84BaLqCzvDr5oP7JWzFX
Cm9cqORMtlVl/XcpGkzP5aOo/o2HaSAKmsiViPfs4XJrw35jjYGR/2vMiJXmQ6ax8zcJsIgMBBRF
6Sk0chVRdevx0Vz93l/3BjtDuRVlvxQHq4ToTSti47WlhNyjbcZgQvO7qSJA/Xvg4et1VNsK1/sP
NCiQJmwxjfGEk4SznLrwW9e0ZubLtLTz+ZnEgtih/xeY7BZyWPbGPxFFPZ/19Gy7ixkYEY0wDk0h
t675R7n6BvRIpwRhfmyuIDJU5+Yfp9ZHMQ84cnMasyNsoIqgae9N0Thc6KhYGGiBWs/CzkgRk4lp
ior9/umY6b5gygiMf7AVhvenZpatwSkUOs+67SeQsZz2fDJ50tK5FpQyIXu4OZdj8RoqzIhteGuT
/lp4PI5BWNC+Il68m06LZWE+mALwqhZ/IQIFMuvbERGYEx6gUl3I5jWtzDPtgZp5h9fAuG4UVEZv
SCNcu7Vufsgb9mCMPTG5PNSCg1YIAoxtiYO4iyHVVpjuObQkJgqxXHQBl6G928IUUFzZNQqGq6Mi
pkeQGf5/mZGWGAyc9BwimC593n73gMcmvO481RzKAw0CLZaLHA90GS/YaJjv3+bgUyJlRjVeL/q2
/vuXOxXoIUOD3wRz2Xyi3LIwUpwmUz09afOKfbqEaWk4AYlzUjSMEZEKy0Ckc0sQm83ESd05zm33
FynrzrJdjsHjFKXrnzDd6JWKWsnlcSMUTa4q+uup3sT7uKDcd/4PDDQy6ROngKCOdO2TDU9c/oyw
EwhabmbcZA82By0+lRIEUrtwqyPltqjbl22GBnxyyDzUTDwJO2w52oOEtHTEQ0zLWtBxDrp7jOGL
YaNLm24McS9gSb6emS1L9fTlC+3WWenFTN6Pr3KChSTNQ8OpQ79JIdt+1Jxd3sZ6NDf16m52HyCL
wgPO/CW7W+kLNUQrXOwW7yPcCpzqsjRKBFRU6t7zV9Yjc5BxlfSIYLjTSe0xklpBLL1OZypEwKCi
fA679LyrVuJy1R4oVnVEBnf3WJ82piDCIPen/sjQ3iFfGPzcPWSOck0kMZfNjw6LJNt9xP2QEFGA
/y3bebeeit6ERl1ci+9JQWThiOjK4ws5vTuBgTmegK9zhDyE9zJqSttrJZiBybtxhYFjzGbzUzi2
X/xQQMm53emu7Rs4v2ov9MfrzFv4OHPxS5nmjwXv7HWV0ksa0IE7rK3K9Zpj85XInaGdJFcDetEb
5Ak6QvUv42rSG9+SR8FFVPjiiTdtk0bWq1DcAhCZjWPj/k78fIDQmdbuSHpD1WpzwxdpbxiTsoCf
wj2t8+hPJN3YCUJFhRGO5qPgtmdossQAuX9P+Amliu5KOMTP8gENbuQb3tEktI8g+liWVkMd0Tbo
YnybfxHya6ljf9jAXsTk/Q/WSR1hTA9AR00r2pp16Cza8/Dwa5MupKSzKthmkx4Kwrh2M5txBIx6
B0lObGyoskXhmpcZITXypuAHwVgWk0MMKg5G3p9YTG5D8q52sPDYoGCaP6wPXIZ0Ox9c6t8e/h47
cFQt2DHBOD8VPrXMKGshF8D4+7IG++EH6TpQ4a08xPaiR7RtucJhK+sVCw+owFs0yT3ipaRaw1Xc
GjU/Fxtw3eFTCeOSfvojoZIQ1qeYnWxMDqTDJMrbSBaqusurfmh5UA8elLHAQiy3OvzqEtTqMcid
RH0hB1mE5RUqw48ajg9Y/TdpKO06cTwCzaQzUHA6+WfB3Ke+Kj4nl/1fFKg8cWmylXJAKlLZc2oE
QX5xS6k8R0Yf1oYc0VPUJ+eJc3sIVu+fl8llonLeSC4NUPKDzj+r9kYk4uEULFy4fOTLEOpsXzTy
ZfleHMdWQdr8y6kMVzZREAxQ1kHYzQN0e5auxisQ3ijJ+RZqKss5EZmbaCyz+HuM+wWNxGgncFhZ
XWiKRFU1ml+I3sGK9nnustJlOePwg4ssQnAv/BFECcFoIE/jYRVQP+fDer5P3QIPlh87XLmhbLfq
Oaapweg6yMo1oGl3AxE5dIeq2m8FWneg0xT9TVPIq1fWASQLX3OndWUqpv2ICfiV18+XEYYtvqHH
avndLNA2K98u6qWgwK4IguNVuRqPU94luWVLX+vf41A20JAhUxBMkrPVAkn32QjNPPFxwfqqINWk
QHQpZejOxe4k0exIVEMAgQZ0sU0IojLO8A1emLj3y18owc9WTYu6Wn+VODPmb0QBdRsSKaRLJwk6
1t14fvjbLmwybbdCGPzj4jNoUKCGcdTjzkt/WzFNqC0ZuxRkN69t5M8tPBvPHQI9eM/682tqm5jN
7dXh6vd2KFVb6BN7NDQz7WLutl3BgaUFV3TQ5HVLIoViehFqkUUtFQocc3QJ9wIHYDWMGG0OqN5g
kWp7u3f0POIXsH01ksE8I9Vz+6mJLjOut4PkggapuU6Gm6Ffox228m0dEJF6Fcm0Lb2PFbHPDlbO
unpTySrQEnnuFtuVu9HUheSjSsMj880vFSQPCC2LLm7esjUjbo3jMacG60wFXSPEV3DtFn8EICe4
ZEE+sRAV5bTLPv/8v+LqXEhidPyQmIQRjvEckabzkRPk+o3T6KNvf5+fpEMJ66/86ITpIHTfzem6
hacd65+pw3QCQPEOZ8oWG3GOQPm/bjY7SOdn4Q+I1eDnP4TzKKLLTHVP8OWSNkuXria7ahI0J33R
av7wQICjQb+JWPPxxzGn9Yieh9xjKy5UjShCEgOiJZnINeZih2rT2qKzeZj2i+BEqoqx65Zl/VQh
YKAVUWcRZr3GhgxY8tAB5m+0BSatNlqFEBi5lrLynm0NFgdeALogRLN/TM7yN8PPVrOKTxOF8Fn6
Ar3MHEtx1RCZmUrDadu/hhtQ/WQsGpHP90DfItUi9Kd4jE/ICM6g7fzEpm/6QhUKcjTQ8/2/sp4S
QVmIQNuq79yacYfs8TU5OwC6N5SPcKkdEcYcrg2My3KmmR6tDvzpNetzEaSie+dvgvyFJV6B+J+U
3lj+uUTdb23eLV9J3moE4VMnRGydfanuBJQihpRi8DudAg7hOg18/XezERnyaYS3/qQ/iYQ8SNbI
UMs0wI5jSHyLlOiU+Ynh1TkKBOuzrPJjDf+N1bRE1m6Z5yF0u0VRMXUVM9++JYUTD4Sd8azT6Y2G
I2v5k983O44G5uSfVmL2o1qWXSN+jygbjA4D2ThSu/69ThefqN877hfnj6MGlAYix+ny8z4EvUmX
ORqjIw1rUpqXeH57tGAT/OaT0BgLWGPQuzlWFGRBGeZdfmJP3TOU7zRFA540T+mp4eiEvoUQLo1v
aw7JO0go7DdHT81n2ynEHnna+kWqU9W3dabmlaMLr6MgZotpRIHTYj/a/SITlDIP7w5ouSRvQrIL
OOAnUG78hZvyHiGP/nKf2yp7y0yZlAptsGjr2s6e1eqsvqoLRNZtp7ENy2mL294e6ej5JMpiIMDp
xwKWan3FToYhuBHtinVRQC7apWo9GIq+x0Y/0GcgV9HX4tbspxpbKuQeiVMh6LrAW+74ziyOuQfM
S99kVCaGLJ/+Gk8tdUAYEfspSyNSyME6xhGKpJMgfWeRO34dn5YWSuci4v07ScW+FTruUL7pMCDz
sbWuMXtLnyJrXr1plKwuFzvSFRui8jNvVOpZ6xqht9iZ/zW1n2BD7IJxov+z4a8rppXd50wca82S
cgPQV/e49j+ynGHS7ji/xdDrbOkVemlxXtupuUmNzsc1lCuwxjdxlk0MzQ6Y6wszry0wXH3WEnpq
Dnd9LzW/HuZf1rqzVh/oETyXLiAjoZteFzs/2u1CNTmoMr/M1BeP5MbVzRXJV0f7Ed55Hsq2mRgv
DJkmYGwwZ0P4f44zf4CJJQC5b0Q86dDqZ3FjdbgZChsotx50xcnwu1zVIz9Z6aHqyMttRUSwj5KM
7myoIyuS+afBjV81Z4MzHWoDGlcxQwpkS+WHQRZTAr4/tSVdcujNdwDTix+FEIkAhdecaYribLOF
ggSuZpdctqxXkJwoqNGgdxTAM3pVpcu2m2FhlXbSuL9fUX273uR/YsUyz2i7htKg77fKjEn1tG+P
s7A6TpSsNszeTlN4zXtqG9oHWfeErFB33IRkvOYiAacSkm/aXU+lZcmuZRQFcH9iydM0rug2ZCrj
Lg6ZFmv1jaN4JnCZknpTk2ujIXGvYf1hFXQCLbXBkMeMwhyzYQl3iFeLxfFZXqL3M+gvxnqtKSYf
sPz5ib+VFqv0qB10xH53ar8nrH9kNLDNKvTQFcNTk/Uc4wj0AcYUrs+STIcnuu8m/lT28lCpzXvh
7jPhZnvBWYmWuDRYqyMMJlY6PUMm3H9RaCpMhueh3B1AbaZ0tB7W1AOgTL+G9JSnl7cWuuH5LXil
ifrpcjdPYNTFuJDke0q1KZskjOsb8qvmGRhhWPONITgRgKXsOtfAiMmEP+Es7phk3N6z2TQ4ksqs
ktUo/2w8Cc9BqP2r3qfncAi+L17y/WwnvZ2HA1HG6wo/VjlkRGHTB2RZ1X6XFzN+T76vDOt7uB6a
SjqkhgDzBekEF+6hYhqt5br4rDr1bKDCjx8T5uYBlYDgzYbafpvTl9wmjgRq7tdeXRxmGpPJgrKM
7uGY+hKEkuZn5EJ6bMReBP0rO4bNRq4CYK2Da6jL0HJCTFA43b9q7kP8bmTBJhcJJyDtX3uOy55K
NVaAsGfjSjFilxwpODsQyAe0GoLVLYBhZ0gmDn3CxbWqITgpLBNQW/019Ao84pXyMsna+bkYAZ30
xW9vNr/wMdff/fb5GrJmWZkJwJJjtJNVKZWlSsXaSJvl3QFF56KyTl7n1WJVz9lMfReYRWoWhv1q
PxRO6/jGVVaAbJsvF2dicFrgsgM0yXOByIt4AdRp5kd9Hx9vWaMFn6cukNbG7IElA3HZ2FqA6I+C
bhfr3nUsvpK7mFTmNhYf1+zEks4yKew/M0o1xd/E2FXXSCExhtEOLl0+VILfF0cLMlweziRO7WLN
qEcp9g4g1UF1LhFL//TdIlbcXwxqIq5xPVnenANSlhaNydoB2YmrwBOAdhrnU2G2g4l9wFiAe0Uw
AYKxY4MMRpa4fiac2Nomyxk/PAyEZc6/1GHzGwN6kwXyGLXBXdf5zjPf8YfvkbuhiJJCSVcwWFAD
chFEw5XWGpvCj9d/zKWOA86yWO5yhleHM1qZKpWE4+k8bQXv6XrtkhnyWevF9wqPkC0oT8Xr0JoR
1aizeXF5358CoM7NHozEBvkhQyJ71JhedxwsixFlbWBtHUeZV1bn855JbogCZAJ8IetgsOsnc4+O
6hh0h91nFgNEFAdqiCdqw5wjn1E0i4las2ey0D2g5ce27T08wrJVfMYQj85/qN/HaEvjVtdsFm4w
ayilcb5M02bCh9NFWGuQofMwTyCngG89MjH9Oq2mSmkSsxOlUV+pjE7pe1T5YjN/K9KVhV2e8dGY
olZBAyAyN1vJdaAA6UsK+uB1aD8V9EvPqFi7ifjNC54wHfCeKKQgLUI1nUClTEDQeCROUeEEZFTk
YnpnwusYV72pRMht7GerP6IpVJfTfw9Sjy64UqNilhRfMIzL/1h+N9OJsVgsSb9WJLexvmmqAJh5
otB6v/a9w6jzb1wgUe+nBgy4+1c4tAXVY3rwJs9MCsNaPXaLc15qhpG5foMLNE3TtoQQMtb4Ez0Z
7cwJIjSXst+1b+qU6z4RtHUfHNA5gnqf+7CLDVlloUSKaSgZkjdLXFcN5od26e3BrxQPoic63Xxu
ZcCXuTAP8csK6j8MiOtix+u1D4nc4nE72/CmyQqrlikfc3HUoJw7B/tPuFNAnUjxS0HR1cNvZ3db
GsDzCyF3L5hR0Ukigv52t9kseLi6WaO08b8zSSLvg0cHHxwKzWSMehkaTQ2WMpPolDCHZ5nCZidg
8gTN3jT+AyZo/xgjrxC6nE3UVdmQROSHUUIAPd7L1TIVqWU10pHdqQjwt1uS/gI9ZRapEVQtzKQI
0DAwliBspRbPMgnka+u1+bOYxvtlQoqaedEsXnlRmFaRkjdFcgycrOnZ+xd+jdrso/+LfBI3OZHb
yRCaRyNiMnng+GpK92XTQDKYmrHXBpzWwamgw86hNwrG+E3W3IeSi2bN+TFMpAqccX/NKG71m39x
1H0Vuair3T0aZ9qZInFlkW3n4yxpReUM8KPQi0nqIsz6kEXn8QPQBLWewiMRgTWBhEbfM4wPKe/2
Rf+gt4AeT7ET0fSIS/J9imhHc7hXP9RUdCfvepNubS4YXT5nAKEYvq9ms/mC6pf02uI0RtCbV1Kr
Xo6czYj87S8ZNrPyON3plWs8anUHGwKPe3haV2CMOCm7BodNsTKYAgBH3TnvhsEqkhFmHaz9V0zp
1EIzEdOGJQ+3IBnahcVFGO/fe8LSOMnXAYBWI+txjHXdtX1OFlsJdKU/OvK+S+MURzLJIaTHwCyK
3JPrs8e/wB/O5MJ6LmYUDHMgSl3ify5zEJvkdQpU1YOig/0mbo/nBeT69ejR3pf/N3cCcTyToG/W
dIxxW5sOI5ZcklcewBgD0+QZLiWuHfWzTstRNUil8ud5pBjAckzFE6iITRALVs+f0sVEfvrHC4Dr
2lyd7IVWyxI6ib96ZfUxJPjSOoU/5RV5BIdTGMThJfnJT6CO9fGfZP4XNWdbd5yDszcHkU9czcZt
IrvjLVOG7q4h4mImsFOhGWHx7sR67OsixDoebFkhN6zhdkNJNJSbbRz8B1KtEeDSjh433vElepum
c3hBvidagXB5NZHpoWlw1TriccCfnjkLbQIaWSo25+IIdqpMoAHiUHu/YNcXUjY6GBN2LwTJ7gLL
CD/zLjdHrvgVtYxwCP0jLpbD5syHlEolmWwI33M5OxY7e4pKn7/AgE+UcXAehgajh8R+9oSDp+7M
mc6qLNuDOoZrdFIWBa3jgrT9TGnsgLltNGXKdsjX/t/vKiki94lhKteMlVn/uVeu9WyKorJoCnFK
637dLtMs3cT+q6EeJnKQZ8WoKrz4/+EZLg3f3lED/7y7pRZIGkEMo6siKlnB9XQTvGsJBpYcMDcw
AP4RaHVDISiME3ktJ4/gTKEaAMki1Np6mZXgzLPSdjAJZEsbJ8VG5OvznTlUIQgMnSeizkqh4cHj
zAjkDMXyw6lgxEsXwGJi0mWXVNkxG7GORuOpOb1zmIkdAT/l1DGM0fawnXY0eE6KKs906KC70mJ+
SOXz+WyV/phkg6cMU01iUnj4GYz+cuj+TsuSTgcfSyZd6gEf1jJodhcDxxh/2CZfKTuKIhMIN9uR
zhlo1zrTjyikhEh7JJ0wvUyrsLUr+Ca8ZXaseoF8Nmq9ZYmkhwcas1w3XPPsj9sJjvaOPidBkn0T
5nwfcHrDQXUHuMPHeLjqJrXxutjDdf+qrhvp8uy0G+adq1wx5QI+LRaLoxgMVhDhlRLaeIJUqHfM
DcBYM2vZekdhQWizog3oVv6ZcA2EItInlOa6ih9EsiL/sV4yE4UYj4fCxMINimmz9bFHtgKk1NgB
rYHB2nimBNn4WiZQ3Xca/1UDjKMoPPjaO2L8d7YtMbtaM30O1Esdd3udh04HdIGKerrUhUWO6h7i
4+gAitpKsO7yCRvKaA6sKdjUdQvsjcoLq4PStaymSSC8kofWFcvipeg5n9mVZaMD0p9Pun65sF58
2q8oxt0PYuFNM6nR7/l/zLINUJLzPq8yCrNh9LHv70orGGniOwXU9f1JYj6YkcXe5+mu7A4TKWhn
2e4PgyIx8Z5AuQL6CaQWUCReRQs8YLw7zPkdO45ToL2EUsZ22aJKFejmhEw/94CpslrmbwrGAIF+
+bwQZrfonKtaI/3SlLHJsGt/u397QcHf37NnA+PgvEdiLaVf9gOUs0nuERhJD7dMVjjCcsONwXMZ
W2nMxo7Jjb9BAq1m+PR4aR56EZ0lv2kB5f/nnrIa1sWwdb0EO4CGILWpO4p8ivF8Gv3uMEVkdIE0
04yRb1iEWc0SCWbnrjf8RlI0R4DkDYmPv6KLDNf9MccFb6wZo90Hp2SUnnXeLAgR1m5WIcXPUspk
7UQC6kF1BfFz+SfV0YBql/W/5xBpr0kYh7k/JfKAF8YDMXQbCDrAoPybxSU9sHSLy6ZwD8Rye2fO
x47dc8tLvsWuixxAGnh1XfeTuq/8No0m3HZqmzznVmJE47ED+FITgTBw/v3gDhBjHegAfTs1cnyO
eTCLVLznUBWiEDYWBNGOIYRavheAoav+r49CIvyVxwadHihzwPWk/371BKouW0L2cgocP+r9HWpR
0bgva4eQMddpPtQKyWeWQvUies0OvYp9UBDv9QHypI1I2+Ne90O1ygUWscPiO0aVtcZ7IQ7ZdERJ
8Sh+rWUYXEYZP0CDzgMGmJc/s0Cghl1h4KWo1sB6SqXmU12CnvSZx2sQOjx12J/iT3+rrj4gy/wS
rQ44sUn/eCm2Yhd7eSBR8p/us/wITTlAWU5Md63x0Od1dqiz2PQoEyzU9Yj1I3OxJJAa72lwY9H3
h4Epb7hDaijZVHdBvYJ4uZ29KArM1ZjsbazV+iSQTSOdz1wxVpo5q2/OjJUCR7oNrKcbxYhD8Mzb
9KkZ//LLi+RpRsv2VBRG/uMjYbNWg83s7C4ygohESfu/IN+vB+8FbcFPYnK73+HBJeDnzuzBAPNX
4Uh8iTJJZa1dqW/+wfAUqp9noR79y3rbmFO1VZ2OPtwW8mLpdBvpdXfwm+bpIKv1+TKCGPySmuwN
qNPvUVsmGrpn4duSEc+41ibYIBguIlLSUCe5PnS5Awsq7/sJ7QxCTFb8zihgdcc22mjeXtpNzE6C
CUyMFXXnP5cuY6blXk5IQT1QRtBEFQMdty+XTuoGHfaQpb7PGWAKUQXjL7jLQu6K2d1wYplxTc3o
IHOdrghI5wiwHzXoiaEeLnh09roYRaLmdfGgd9FhBjOQ800KaXYiJC2ScU4Ezv9zcI7wp05iZBjf
xdkUiDMqhZ7xk8u6SgapKziVBZmdeE9tJZy5xH1dSOl0yvgoXrxt+Sn4IkoAUb/cpNAeXPqSoq8c
15cseZvYFt8dtQ+YaxAIruf3Ro52jm+1dWbpSfOyuzxjsD/ixHDAknIadTYDNgjq34Rx7R7SBGxB
S7lQhJlHO3cy44VvXQcH1c9VTIYiwPtb4s2K6r5F0UbfcCMW808lu57IpyPMp9FIySCha5T6bRbx
CO4uS5xmMm4hCSaISN+9POnzp+fMh9JU0iY+jcn9qOGq75WStjHT/QT1KntKXZtrABBG5e0m9qwd
K8GILzQS+WMA9QnSyEgW+t24g5qXmgh2iwmT3BfNMZSbtzTzTlWu0DEf2hUyrwqB3Fwgv7BmXRNx
J79z0GvyLQQ+0OCgtCCm+2NrfikVauC/raBMbZpvR9ZSKPR0Zqanq8/XxBJEDx71BYDMhCCD93ky
mS5GG37g7/xpQjDVbzSJ7tk6Sdb5syS2Ttit6SCM7g4K66YqZosWMdlovZbQ9TznugRbKu4W5mf6
wYv4O5i5/R7QqQpfZtaWWIPEPz/fxyrvcOq7sgdN4O5lC46cBVOSophx3ABRaK1cscGQ2Y/IrLYn
bv39vgUddAfV50RKLiLQu9tGtVRygfwSIkRM2nwotfKBFyN/C5BrSM8oVwY/CUHIBoP9CWyCEKjI
unJY7l16bCv5UyM/DWmYAl/QPTjp65UiyZjMi83HO7pVzUaB3zIbWFml2+6hKiKwSUNKwn+CXmJg
TnTLLoX/85gze72EQd+YrURpU2gVRe3YZl9ectufElr9AmxORS0gujmTWnVoiWDD9XhrTK2taIGG
dEEz8Oq3ljJn7RDftpCE0fX5PJxZk8YelAPFI9fe8V9+gOnpnoMXOMp1/e5hmM8EPr/HLUMKkWNh
R4T+huQ+Ny7i70vxWAmbpxBuYRtVH1woTnS6QjWi1JktFuJMxwQi54g+HIjbdRyh2Jdt8WTDYUIR
jC0d9q62xIvvROBuvVSeKImkiDjwOVLu+9HhB3Iq4fA30+XitZNGiH9sSMbtlQOqkxQPqDrl2O2T
wp51+KYPuHeQjid0yAQCcjnLO96CqIBIY2L8alt6MJXK7TEDGgzodUnpRbQ4PHOJMWupGhdwzncV
D4ZROEvAOoBEAgUDD46eUk7yMWnCdXLOWRqQOAU1Bs6tfCLsU3PIPBCFcw6GnsuGEnFqArJHEeQc
KXNT1xgmeoDG3j6ISR9/tz6/ZIhCoLxg95mfveoc/4UNE9gFVQQ99twSgEUrFQvtzKBb2u6hIrfL
1uOMG1wz/wTGZCESBS2mBm88lzIAUrpmyCUg5CxDryAHBleVvgyMU+/XUzG5ytJK245EpkFMC4y1
H76enrGqTtAzWn+yl/9DUqUdKHUf723R4sTZXRIdhGHbw9Jfvm1O0OGBR0rIE0GHpxpjBSR1YmJI
aMzMLlFSAhkfeaEN7RdjssBRQORbts0yR0KalQWCa2A6JqJ9rBex7zfukN0IwZQ96LeFjx62WHmr
X9gQ9RwQpY9L2WLLlBi55/a7X4ZWSdAXfbAxCtWTnbqhUIgkUhNKYYUpyjbIqzWDEL+0AftnFbhG
Asg0sm79BTPgDBiYCQ5jgw4HdWpo6OOw1iXaEPzd2mp6DpCIEk9PmM0iK6lIdVgIJoiZDyx5FLV0
NVh8jZAJuJ14C7ZxHtUmvKce6lfKfgbftNHck1CWPId0IM8k+t8Gad2yPKCFQjmctBNa6pPhWB97
hDnTpGRgsudadY2CkWE+aZLr/zLaFKdhbK0O/+TvpMH/jmx7Lk2kfwhQOwJLK0jDROB9YxF0Vhae
w9LxcP/VwWoDEB4tbmZYDI2d9xnqSch7Z2xpCRWli2wkmt7NI6qfLoQAyMy2vsZZ/0YHM+nar59N
NWDogQPLaZg9IVRN8lwaK16HHZeOAhL7AslTjoR67kZZyeQNw7UL+u3fgVESQbNJn20qB85UQbtE
t+CeHsh5Nwm/g9KREfSK0uMrK0Z3Gf8EEESUqUsZVA25firjdN15h1Qb699e+kx04goR8K/NbcBO
Nhl5Gc0jjJR/OywaPW962kvfvQetrue+lnYgRJ9MGUbi1nrjOC2xFs5Ve3Vrf7UCtwBhP6VznMeh
DhNrL5UOlLw7UyhpkUt7NiNWUhv9bJhho1iSHkpz8hotsyK9jOiEv14IvEaBwmlkMgqAUkyHfrjj
x2RzWKbCr7DUZbTYAARIbGxOexf+xdg2ZdWp6ijr1OlE5PThpIAd8FRsdfRlolfMRiqAiDqKN83n
+GMB2PHv0GWvleQg17potirb6aKmEiV5peBiJDahpCHQiMUSCTgMMKNLd/EbXcAwYyKvyE2A/5b9
uUHN45bG7a2Ixd4RhYgGJQU3K/A0kuCpmM1Rz4bT/bHmP9nnHTSVMKqnKKTHdqSMmuPt/j5EFzyR
qAeKqJCNitrNdoD2o6U+/95owsYMy/dF4qEnuNA2okiQWshiTaRdGV3zaqUI4OKi9dtr5B/P/MEY
xfSkvS7IQbgAuD+kRRKyBrcwkXl0kY5mQoQLHojxrJGaFSsgSyu/GexKo6lkrdWbcNyd1lnOpQK3
vaKrJX8SNEVGoCI4fs6EOuzgyaezgwViLq6OdZJgFtMjJRfcTLr5SwmKHZX+tgtXFgg9ElwoH/ae
hNFTQX72ha+xoGYJ9rTwY5OdPtXXzNnFSp8fMHh2LpFUvpk0HXlOTIms85eYTQv+t7r/U+vfBuNU
vij7cYhSo5fpdIG5ylXUOMDDzG110bSIoDBvb6Cqa+lxROu3qd+6+9VnuRU5C22pu/vZSglc1QMy
LdH33Ww4TtKOGsQkoLn69aos3jbGkykc/39OXX6EmMorAH3XQFe8QJMnw7EUkuduaovEELTDhiHH
KIPWMSWXuQ54oKzN0BYuPZCvWTFHKl2hlsqZClB7TvEJLdSmQjS0qosdP81GbeftV+L/x69dN9ls
vpFMTNmP1Xe1mKFTD+w8NJFyHbr+3WXCarIpIDa5BPHetGoYyaZgeqnZKWn9AyrTCMojULyZhs6V
6rLKYUQkC87Fmb9CDs07YJugLWs9gw6jBvGo8ztm6EK8OCZqmY3AXFEa+aW9rBZjuJ1FLytbEViJ
dE25FsmlsezS6hMh9EhhNogGKra5w3NT/C6b2QoKaCY/avihbJZv5RTNCEdmMutmCYA0ZO2fiQ/H
yksnUYVN3RDaDD5CCJKMN1wa+YzidX4Zr++wtqdXDWyaVjxC1iSU4T4o0nqGmp6GTNVm38g55CDD
j/dFbhkyuSJebUD5CV4jBmL1/FX2K09ZYhcZycvi5hfFLoVp2HpGOOsGZvTolzAXIt67tOYJL+bZ
csipNnr/NR2+A6PjsxC9ULMKNBXKCp1wsdr1M7WulcZL3wJzuNEhabxqMvcyo05XbuFO2kxLFnXP
h3NsKoDlYiNHOdBUYkni9/mO+Fl0xw86cPmL1LsBz2p5bzGAfQQCUQf8uDsR0mDQ7I5pxAECylSk
ceWjgi4T/ij1YtvOgN7n8u7L8/LVaq0xi1YPCZaF9m3hd+HtMJDClT7gMakA/chSCmy5MC+ssUcW
11t0gPulxoT9bO/2ZPxvrwbzyg/P2bz/hImRxwIXczBOZx+4KqEQgruO/oi8/TXgnUBK1mvoUhzP
aK3VP4h9LiZ9JuDFvr8Y67NazPn9XgKJCZLTJYCV6RAJOPbtpYoiIQ0oDVGLaFTWXIJ25kKYFCQ9
49uKmdNuE9XlFeWcS6+NHSDKezrX0hHnY6Epo1LVtssFqDZm40bLeB8pQmvoL19h7uUUMuSTxxPq
7iP+jDik7XM50tpGm3YHhaZyZCoX/X51cAI/vNE3rIcWMGPlsHN1CN72OzNcVc75u7a0bptPADV8
gYyoP5WjJrG4Nh05YytajSBkWiinUaRSS9A9E6kcDCeS/BrIG52Mz/YuiqJaA1U4TaaZ3p5xtKId
Miw1sOhtjg9Wa3NLDIUjSQUYWwv8Q5Y/mrf5pDcZHxGiwCiTwJYPBCqUi2TRd7V2z8Ws0u/+7fng
JAgR9XbYhEopkQmIFHZGxyIf3HFXBQLTm+Gu94KvegS9fT3BGIpkT37rAekl7eB4QFTSuSjesb1v
tsYUbaxrrRKkAZ1mT7IWQCEsJ1kWPRKm3aE/WHiGCq4iHvAN1tV9nGBTRo7AxOmkZFVyY+ujXb06
S+atIXe0KHBhsQ12ou5wlmeVtgQLOqYBgrqEngAIElMp/yQ8g7+xrAsIRocmxQsBQGTs5i1wtcB1
ZyW/gavnfdQrPipC1fW5EJx5GeRx4b57Iv1sJEY3yCNtegnM8HLBnuBzq2dWqveepioECJq0wKvR
F/WAzXGQq+3Cz8Sk5abiwpNSD66QcWKVLDj7MmduworMKqWPtrZaVaKvW120Tq6inHcWXhKcD0oI
UM9u3VkXJlgCMZyZVwbVphDRRD5sdNOvkme5TptVFRDrfXA1ocvthqFkwlw8pCMpUUKYhdLfa/Jt
6Dg3Pca10I6aMUZ/tt5SwVKInJf3MdZAKeDsYnX+mcVNSMIf890pava3Q3oD+JuBtDqrX6WVgloK
uLVd6fBNsq7TZdapuqHd3hlPPoCmLtWDKCcHkJNqO2bm1Fsvfbg7xduSEk4ugmrtKV685PGOHgY4
5uOZEyfI1rVp6f7yH06RG/IDZt1BUU2fdynIMXUBG7c8DyheRff23z6KyfbyWNbDw6dY5XeKiuUh
x9SpHViqUo0IkoMA3+dTU13Abpk29kjc1dYR72oqDuL4N/g2zT4O/ssnQDAe4Co8QvzPX7S4Qzwl
cBjEMCPAdqtMvu5O40Q13DQcIQ3bJzKjhviOoP9T3vJsc1Y2uCb49HvMcf92O3V/NLJBRjR+WDwE
cyIOPXqARiikbV2irrZVWn5E2jEqyqBEBb2b4M45A5hINcg4E92BIUgHgPpTtpUQHEaTIaS4h/Do
iRJLA5APo7m9njDVYoh3fNtHMKKv+xvwAASuCiZxbmwtvRH0a2C4fLE2iUKm8WGcFOaFxcyZCQ8/
AZtGdD7uUsVjiEUqBfSif1DrME/vLLtxU4gpSH9tk7R30p7F+zwkbVHHYipE9/XQ3HMS3kdWGyAu
1Bo04JVj8IyN3SsRBlaOgn11BoxYjiCxe9ks4mP9GXkXy4M+7AqWubSPBv3TP+DW3wyntLtCx6yq
aRjvD2y9q7wM1OVycbHJFvkNP3ACfqJK8Nm7O4Sem/k5qcZtwhvLrwQAx9h5Nis3wIhieXey6RRo
noVdqugUIN0Ofsn8MlrPjNb0NZv8dVnx35FXEbpUYZ8o3aD1Q1ZBkp/qx8S8eWtGF4LHr0P3v5xY
c/aaa9luAjFamslTMZoSD+z3bxS3QTCpeIRwfkIBqd6ldz9J0qQM3rcHFCrOcnWyOT88K7GuWrHI
trkNwW1PY9vvoWGvgF0ljQdutH2tJhpZupD327w8vO3RCB/CbqLbbi6AT8imUI5BYwn8R5AbmEPX
HTdjjAULDhpEhZ01Q7ZIH1OM5deYBps+KIMIRcOIFxmhKmz3G6Ggg+4tSKIzrEIeL9gUhdqTemUx
ZiEEgXKstJu7ey/P+iEi0aIv93LUIzIEy3UAVLZ+31jLUn/Fytrdnja8W+JzMNpRI/OvmCeGM74U
0PgMByNpBDd2mkLNas9n+HuXhKj58nxOOdjXe5n/igfMf1uGsskM2WoPEQAH2tlBgC7uRu4Uezr/
M2V7+oemH/mavavIpDILqZvVx3xFAbADKXbwlZ2hC2/1x2SdRxUC/00Wdaup5JKGJCuBNYJEVqNf
NcxDo3koOQxLkY1g1H8wrHtMc24V/SvdfwbFX40KlXyf4gh8n+RL+Djsu4P4Mf38Nd1DIzVvfzyM
T9uD8zLow2z4KED5h6767ctnCdjVo1yeYI4LMJ2eKjARZTu4WLb5lDmcoTOyh8/HoFqdr3PRXFpn
soQb/JXc053rSbkLgg+mv/zukLkSAJ2/9m/0qVpAqbh41g1QE/TLYPmP3AnZKrE8GwACyTzWxYSq
ZrxxyJDSfDtTo9AvtPxwoMWZGc2uVu5D05k6BjUujc5FNI6L3CVXni0rPJpjUxAi78/aDNQrgCXR
cO3cKrk8+y3u/BKwLFzSqxzYvJY76ZgKv1/xTrcxL/rNEg+aJWTn+9MPKL9E1DxNTr/3eRneTyNx
l6Gqmf4PQCSNWTg0YwF5U9/NwDfkWdLIsvklaOVYPILA3QrAdcr7zVwUUwT1Z9T3HcBMdJWCSu/t
Mfc/pQpbrK+GcyrC7ZmzEUVm2M6RCU4nrdPO3VdsXgsPVfbukLDX5QSS7ROCU3psusx5bQGwT5fP
4ZSKVf44hRblQFspYas6HKvi3rtY6KpnCkYs82womTujwYj/nt6xtmp8KZ0JYxgZLVB/PZ+8YqII
ueVmLqotHeXaD2pGGqOiY3yaYQN4VVIF6iAemq0X36pzeHc2NUkev7sSbatOSdZHO82eY4LpMELS
m77BQjCR48uwWzgC0EeZx/kFqUip6241Wqildm2Iuk5LOvFXbHTuNTZQ2TYt5sRZXoSFHAU8H2g/
yfWywdmXC57MYCzFf884f08L8pwgiqD9rqZTDqST+2iWyYghRmocMiwslRENp8Li7H7Eylt+g0Fz
2ePh6Mn6nI6NZn2N9dA2Q8v+SbF++BFSkFIE9bY3T61L9oxZEyaLhrR5SNzydw2N5uoEYOXFXRS8
KXrDKHWGVUJJRzehOc/+1uAKHI4O+6P/65C72jlFh0CgkLX86W3pzZ3R1l3iLGLkewHa8wcZg0c7
uvrkCV9sr/j9wddwQ4Yj2eJq1cyTXJ+fCamqkNcew9Gf/BsKT4lO9eQ0P/4MW+3NawYXCxN5grqS
SFk/balrqSLElAzPLyB8Y7I6opPt7hvoxfoI0gj9smq6aOJ6RVO/yBbyuTvuxnm/v9X5pqbEQvNZ
pXKPNWsV8CtuxfHKjiM+SRs5PJ1QfpipgCXXYSGwsYOZJvvYV5SR+1YENk0TWlio4vnW8loQiP9i
8YcJh+6oaDYjFZh/lgRrZS7/IUTYdg/+t9PSWB1vKUe9xYz9wGvIs7/mxxXKWBFG13EPJi/VVhWO
JECxbKyNC/rtCtLztH2Y8ILCz10O5IcRbo9ZzywSB/bOPGamAffwg2+xBIXTIIz133T0EweQ80SL
4sl/BziiuX/SwTHjq/B8LpIdia8OTMQlB4/yZofmsweFiA7lZ/piBwmVSTl0tqcrdWvfoTXbUTm7
G+8oXQRYBC6UrBrIiC0SbEUVYy8M6oTYEUdLo5+kG668DIzArulaaLLpNyQA/+4V508gnU0Egago
UZ9t8pqwry9vCa2T5LZnmqEzzfcxwV14FUsZtQ0JaPwT8YB9d1QXOw+qYZhNHKEs1dbPxG/usxBM
oPLMMbyoyeNkliRGi5K5YNsTqWbjpWm+VjmCv/pIldPe51gr+zooE7/Udvw+1izwNhnk5ceSVN0+
9ApYrstttLtzE2+f9juI1s9KlSDArGbrfg1VbTONm+CS3XwPIfOjXS7Ma1qJh0y0+cMlFjmdkdL7
V/xLncqtwmo0RvJs59eiPqGbLP5EQHajXRqw++YipYm1sa+WH6bKZEzwFlhqLS80jwymrXC7+4pS
b+STPz3U6bOAQj5aIErFv5jxGLjiC44M/oONdBB5dMBNV0mHwmqp7+qNMEV2IGdAF6H3QVBMehWx
A2fyYgg7iP9GPoT6GBLw8eonVED0sGUYPpKNjWH4PFKeYcGoT7Ge+2K3fNTZg6sJdIceHZnSOHd/
k/j46sJZAQ9DchE1KtWlGD2bM8PHFiYyrlSIJ0MbTJjumlmFvMzJ9DJG3yjgN8oaUwbLFaHymIAC
GV4nJrFycQPXsY3dKT0qm7H5o9fDPidlJmATbcqVlP2XIEsT3k1aCantX7RWhtOXlO7abQ1lObA3
ziF8VDsSmastUalm8JIi84gWzNyG9ynLh9sL4MCCDb4DTF57vz/EE/PrQwR5epGi/3gLQjB0eAp+
e7oKG7fNW5zphckl/ydmldF0iuVMay9Y5Aw0a4aQx7VbZFfQ5T48QJF3HIIG+UbC7Im7bCfqgSiD
3SshbZ6TSDgL/aOmZVXx+X4jwE4BMpL+vQar+rLc3tHPs/eL+/m7HS7mS28FcTGI+/qxjMjygz2n
LcSUxdD6+9TFk1ZtCNmqvFMgaSiaZH0Ud3zg7W6pIl8q1D/iVvzpvofoCzSI0qhQwE26vYDiVviQ
kJsW/xlwGGXU4DuDCqvQdA4GWP7lMOnL5F74Nytk210c4lmmbz3ehzSM0Un1/wA7IvUL0grO11dn
v45axVo45sOW7LSfVvcW1kAPWSSi+cOX5sfo0BhGrtFI2q04VkHM4vf2aumVsH29NUv1gWv6WkwV
UWSw2pYzJ5fH5QptIoSMN2JaOEK1EQcWeCm8Nycwvk+c4htcLzlxvueFwurof4T7Hh+Ir54A+vvU
IdoKFgPfuulUcMU8f6u+kiD5BNAvSLpnWFDg77rwkHhVC3+rvoYoqcefwKBV+hVrv6tbTGG5ETge
haTGs7zg/c6Di2PZKEzBFSQA2Ae4yz4W1bH7sU4S5kHYeVaFOlCV+t55eSOEspSSKwo/7gC0eYcu
+DCr5SQvsd9tK6HAfpfaM+muwFlhrUN/PIa4RDKFoePHQbZeSva5gdd/X15zOOup4CqW/1iv/MLt
w07EQt7/s0ZEuVT5dmJNmdJaIls5jGP8sswJfq4lQQdokY2IeC84lJGwIMzI4irGJgIfsfoy5Q3s
C29jfk1V55VCnDUqPMMD5hV2kpNbbRz0JHucarMxwyDNUmn/fZePdEDXPyEM+/7y8KuIg3UMNicR
5kxzWbx/0GUEgaG+62BTe9odVt6LVCNUB2pM30SiLM/zZKzM+N6jjUjLoJpb+eCxUcd+h7gBisul
lSZ+FVEWXIldMjLto+MYGAODmeJf+l/+up28CzusAfgQQYImar/FvhXcOqgxaKRabe5VqYiCGcBb
nysLLYgXBsb73u3cxvU2bxZshQImK1au4q2fAt9TeI8RjOJkc3V9am3aM1GvxJM8hMhOzzM5NUPW
nsGBII/Fmo9rDyiGoTquMmVgMhD1CA1bY/4BDzdmkZicAMsYCEMkxG7uICsWApxVhVa2nBxZkWsc
ma3+T44ELkJSzIIaDzTAmkRmMUdXZz69oJRUZOqSKigjZ+vSjCNf8TRr0/cTRDyIKnyD5TDGUyqp
gCjlePUgC4O/9RE4GUABWWBAGoJh7V1CZPL2XL/snu+qX6a5JnVC33JzOEVEWdfigoZgFsHcBmgX
dqPffNwO9RH9gZBxXfYRBdlqeHpvTru2LZB8l+d+vMgSVB1Y9JTSosvXb9x71CQ10kTOo/0vJPdp
mX5odStpLCzL0e/7it5lKKWEGfgNe6U3M+MKx3SG1PE2FG9p9WdyrhfyMTjzOPWgYMmj00s+Wkb1
nDjV40lGqI9R7kLoJxoGUDN+0EZ5JYTEPI22sLSMOm5NjezeubNoC1VVBlpgM00WFne07jFbF9cO
R4FCADsUwMKXSHmPuPBHvuJ3j1LuwiIa+HDFAXCXjlYzAa5R5ecbUDrJOW7OP3la0uwJRw1/0tYc
k1vwHsCt5XzAKFOVxDmS/37lFDA9jWZDNU64Pn/bSi0AK+urBFvisKSwhQ9t3lWjPslAUhxlnula
uPAYp3uiLeRxluhWXPGQZLK+3W8Z9xk9s4DKsPfuaLL3sacooIxEMDpsZS/Y5fnhSMfrU9IvjWI4
yBNsn2oAgaNlAxncUdERV46k0uwFVHyYp8Ng/S2a3UuPpkd29NpjW664CtW4sKy4lCm87D7TImm/
/b5v4FuTqgOevbq1NPD+DvZQzhjb08YCyb2v4OMhY+22JdPK8X08fRLgHkWfy2SB1vTHkBnl9WA6
CjGSFeFa8Nn5oLY/YKgJ010kb0m6H/3N6tVWZm6dImTpVfcGgYu5dOT2RR3nduxKBKXL4mdxrrEx
xbDkRufPK5vbwNjhTfhIA4BBhmHyVKxIZstW59S3hWb+HCjA2tk+layNF6AMZ4fIWhg+VGoB+G6e
EdEih3pucP4phbZnzdV7Fz0Vgd+7rVyKHOuTUPqVA/p1+vQJL564GLf9UZTQH3dkiD6jfDYefYGs
pzRko/4o3la0kqhgmodce3tsaP7MNRHV6LRLFEFpjW8pE6onDxMBJ/0713mlQyeDGUNl2tpKvr+6
TfTfajwj2/fRGpCcY/3cn6A5Od9iWCQNVa8E3xASmRMgmlyovUx5fnxKnIy8IKThvInMRrwqfRVr
Vrym5OUtzAen5y5yNoT4tH0b+SDBavwBSE9SLrI9pRA5xIVFOocuMqlSAxjCunT/acU2SemeTTLL
g0G0pejNP+ZG1VmbXX5G9CLdlAaeA+KNhlaIH+RRX1WIcGzVRWcPUqHSY8H6cCrQXCAV/2D3ozsa
ycg1lIpmH+Moi9CJRJ1CCm8Y5GG0voJnV5Tz2aSFnOI99k/8Lo+jlhiuYcaH5lyhGB8+K/yILny6
sDOtQUqnE3YoEa5d8jSPCFX3xsHlSuBRDK1cmgvppr+/j6YQJOFE01tSPGEsuTmzMZNp7u9AalgP
WmlVH6ya+pv90YxjqV4YgkdM4UTKK6IaBMs9xCV/wpraCOe3/K6mZL11jY+GupPU7TKI9F76CuJB
qzmIXH1tk17icG6FxIveLT8s4n9xUPX1yjmGhE8w/xzrcuTgAoq2Tj8L54htZyDXH/Sq/C2UWENU
m0VDJzoOtJ/FW125F8+gHV7jY1jHh696eNBVqXt5G3RtKKFTANhurao/RU+fmwOzisqscSRe6opY
LFl3u1yHzAglPQByVrT63hgR+/lESkwinJIMqg3+5shxL1leZzd9+GvJFE2WxFndLdVb9W7VjDCC
16oeLZPl1UxzxfN0ISsFIb8CkYMsBlA5PimRxfdGMxt61PrHi7ZgRqJAlo9UuowEjwz6hywtWyk6
jVzyr7JsntxpGmuBjL5uYrAmAjnTL1n/YQURhTR6iSkPL1WaOyuMymg4pRjlJ/hlOB78AsgtjtcE
jKD0vKBdU6pWfoeDc+SLFI/9/LGf2IXWGIgLqz6bSl4dH0izqELRF1XUcw5hXA4e38n1ajKifSt7
aAFe1/a6w3nWkUMm8apAtYOxQFYnDjE/VXA3eZmQ+6URv8xGDw48S6dN3mIAuRX4qZYrSS45/0VD
RYFqWzor3UM/cEgB/2qid8Vu0bzsvXAq8Tn5+BjSddE1wDr3Ne01mPcoK7gWAbnlzicl1n8kgeKz
Q7JAwHS5I4vo/rCv9J+iDj2MQJUYVV7Al3kLq+Pr9OJPY3NP4xthrzKI/BfqZYirBpxsuNtYmQ6v
cKendNwUEuZUgYzuO1ujLPugZsxKaVEBQ8RybYNcm7TSHfzEdF3YtTfjrUi7TBGz1z/mfx7PF3Sw
s/QUkjJ2H0bnbqxvXJ849b7295c4RcJfUpzdlAPVdTTrXQSqBc7fd2MSX+KuVUxtYpZWS+bl+Fhv
2S2fmu52mSpVQ7VZX/Zjf2+kGQUwnhHq5SW5SG7jpcgDJGQijybtuWmGFvHdNJiF8SvprL8P7O1v
+7pgSiA1EozVQDzz5w8eyPJknkcCfemuDMO7TyLd42Z/hZH1lvTMdhmgx8Nd8RYwELefC/KVTiMa
d8/iHmRaAGIBvR9LVnk3qgDbHqXt/AQQ5LH0JMJ+BMtHxbz6d8ceRDsSzQw8oPlED19QDS2kFd3g
i0Ah86hx/ne0yAbGXBiCyogH6YSTSu6LCsGPJ+lXkmbTuljNgx0m6w03EKZue78t7sstUqIpEoDh
39kcs5tMO06TkGh7zI8Bd4IRyC3C23QhXVDN4/7yPcxTrQXsKh6ugzSiUPOgyJH1QTqw09O6Jirk
7OHySLvxzgmVjdvwaROgOjvXLLUGvoRC3yaxsaV2D/AYapSoNiz+IY7EoU8QajRzxx+qQ5L7uwmf
qSxMAkiYsgWi0PkUjKT/JjRgzeD8zxPWlk+oc7rv5n7FrVGiIvezyqIIV3m1D9oyfXhnQtqKBNEC
yEkV/OHE7hgGBSHqLq2EUpnQaQZVeZUKLBzALG67a8hwoZN9GlTReqJw2VB+3qV6fxdZ/4R3eF+4
ED8R1BJA4LTuurkDF54TQHRLqM6/60+AdAvLIKHOnpNvb43zzedkIFFAp+O48w2ZX9U0Hs60wsYi
AEi2vWXeSbDNjE2XgvnE7q15iY4RtlacwgA7Hrgq4bP8mt05tvIJJ99vfkXAxGmCWdj+6Sb2pTyQ
zr55RkrZojOs4XxfglDeFo/DanxC/Vfc5i10b3u0bgFNvRgVOE9Wv5u8kNBeGlto1Y7X5mrej3NK
Yx6wT6oyl2GeOnI/6iTfacdhWLHY+Xeuhv0i1189NU/jgRI9q3tF4qEI0KrrbbTnBQFCBYkvGfmF
Y6WNsEVbVTI8Wzv3tmm/xL55flzmCAoCFjoRmrAwr2Wx9dHycYwpAFpSFavYgPoFtU636en7C+ma
bkqUaEo7F3kyTJT1lnb++NDd6qLolSmQd1UheevhvmgEJKnrhRVG5eShIhvGOGYcsMtLs3TVNVAm
9pjIC+5OuvKQVTvjLLNIafiqfCQ+8N3BSq47Y+zIvVpW48P5FnJZy1JU5WyZwF6/cB2pH8/RrHQG
68bdUiWFTbqdFAwgWbohmq2Wj4Wj2rvvDSkDH2fpWfmhm5JM4dV4I9ln6M57UFSHmadFo7zDPSwH
nCc3ok3/p34RKAeJrBZmU4n3x9TXZw/F6CA8/odG6SUq0aHAbz91I0QOmzQX+OUZBIneUZEgJ35s
LUOaK1fM9QV5WAR4cqeZCnl4Pdgn9JiPR1BtwmvEQACcDZQawQHz8eGIDBgdFSRy+7baIVHKbu6h
M86DLGXANQ5/Nrr/gTQQY5LYTupZWc04kjbzRi0RdustZ6CBJH50bkyAGEmPEBB5c1gsTbpmnVZ2
QChld71wOrlBJXlZxbsUPiU/WQHd9jzIhlvECXStitdBjtg5AVFfHoyeEtBEvzvaPjscicMS/vlu
qb1dBGXDdq2KAD8Cam5rD8oiCLvazMjkhLXEpigWg4ssa8CINLk6snsiW5GhWH3j479EwMM1Yndv
9vB3yu9yB9Q3FlGgjy+o8jLe7zEUS7QUwtkf0cvvboQu5dgHHb3RX05FiDfipCBXiXlxG+Kc7NRc
DFw/vVunh8mkpsTqDcRwu/qDwTUjQgRUrezSQQb0h2n80Lsqfrzid6VJsgCNVIk7uMdt9+2AqLe4
5DEiUFkZ8u2M2KbJmPLRY+e9X8QmY76mZ/O0ShF+5C4JaK2v7EmcF7jvlWJii2OLLPC2DCfsd5NE
KPb/48XNAY0yyUsGnHR+1qFUW3NhYiRNlIGjip0LGKVx0JPbMsify1rYGAFxjtGTHQuxEWu9Wnoz
WMecq4ZOV62ehqZ6iaKN357po0OV0ph1ngi8XnaxisuzSdkegx011l6o6h98nMG/CT8EkltzJV/B
NVA4HOeCrJeRhL0nk7FEgkkEw+MBU6mzQnxlHyFhT+RHU79nIZt+Z/bjzeOJIFUpRA+Dpr7Wi/K8
a9WviK8S3nvB1QzwEEBeS0owcnX2Z54qU/x7HY7mXO56omVmgzX/uxa2ofdJfog/cpMRdHfPd6yT
TzNVshAxKT5aDpEYP3sOaH2cIy5fhxKGppsh75pcuesi9MD9J7+DptNhsaS1Sp2/A7YsCMO9ybe8
DeHT5/Cp7lIxRbbwQu5D6XzYEB+cqoRoInzS60hAqVupWbjd/sz/Coj7oPXaLZvk896Vmk1cTHQm
NxvkcyFyWmX6If6qrqF07xciKIGNvUKPFQ3s15lhIEtb0EYPkL4IJATJJW52HleYXO/cuuxzC5cl
YaAhmjz+tqCSRgRbAxWyy1m0xG9ByFjzW6MuJHHRzZlnFD8BcpDcc3gcUT+lA5KbjfaD+wgGKOvn
2AygVWt7D5N3VjbNcx7Dw2rsUZCC7fFvVj/p/3EG1yVzrcy58wMjSxIwAyHzYTi1R+R/lm2EJItW
rt8htc2igs2FfPk4KO+gocRU4I7RkscKluxRlKzAo9Se9PGMoAY26rfgYsMbMVr9H0Wmy+I4swJR
hveHIQS32h2b0xuQGXwxC1AEqeq7TsPW696txA8xSQOCD61f90XhMTYSLZoLP/xdGkA+k8+e4zVH
Rh0ToL5FJlg0Ej6f+GQYMG+vc/y2z6qF+2ShubDibzyupW5GsQU+S47AOAnZCs9Ql0XJbhOBhUu0
ctc+lETC7AWiFe0BEyGJ2IwIqW8Bpquct4Kns4DmI6F8tsf+GxsCNSND4PaMfZ6g37aEFT51xEcF
6LQKgQ4rsxCnDKHJyJcfTSzkXzlrTjeWDDym9RHGbrbTMnjLQ+9ouch26cgbE6i0xwnxljY+ct80
g8l7UPyBsMg9PEhmhCqZ9exlNXyUn7Wn3SCQbW8Twzun0979Au5Vz4OjJB+Nc418Zs+cyVzcnrDB
9TdHuc2zkITLjcecqtzIf07EypU+U9ZyInINMhwcADl7cKF0pbCMSR1MPA3ngee89fZ/ziehFzMo
mCAaG7YhitEj4tYM26vq4x0lWNu1oNyBXfGprjq5HL+g5988deJRpJBzktqzevx+zaBHjKU4KVsA
bRzHmbo7hh0dsOU5FjSO/ETvAYfIi+3oE1sgBcoy5S9RjA2AtO5+Ufd7Md7+Dei9RG8LselxxhGI
RahahsDJnzTLvXTk9OZzMQIiEfNNwHRjNJGNSFO3MRN9TsFgmQUsdrxJXLj4BjFxhvCEl4GMWy2c
MWYZE6sgCy5xGcwVcz+rM6JkrtZhvDyGRR2CEpz+XhHgebgKqXQWMIWQPlYBnifdxm1khdYHaKZL
GvtK91SC33YQcY7RQbD/9rPhvfxE7nmA4RwyQ9+joXcM4BUlQBkq4O9KSz9+F3crOAnJ8JNQrkca
8n50ZOjVY/SClWzNmUG5sx70FV0smvOF8yfFugD7TYfpz20kO7vVvC9sf3RPKnoUa2HmXI4+O2pe
kHYyTvoluzZ/s2Jv6Nfek/jOrh1a4l+dm+Kwq0K/xGO/iz5z2iECGaKSrA6b+3xj6PoR8lVc70d+
8qcB0lIF85GxVPWoo2Mu5hy+HFfp++NyCJXOIqEHbZBBiuHN1zQ1xPSGZIgmYsOp2ITe/EAsXxuC
fez4D08oK8OAMHqCymgjSVzui1D4xjHXA6pCWnmGzyX7K977MgEhDef7cSbNclVqMsPEBzOshdEM
AHT4iBC9m67Bgqu21twvfnMtlK3MmtKi2Aeul/7+DdeTq7pP/8UY/C/bA+a8A6qScX58xPL8eKiI
Xh7YNxky8mmz0n8ROI9+3xOiNdT/a6MhgBC7QiJg8pp2wKXdJE/rlhjIQxdnSMM3iVDtpxKWb2y0
/i2ON98ER2JZnwyZXVEw11dWy7KV7lGGF4uNHSFP9RaN8Ce1xo2Uq6+6sWEZ4TU7PjYLl2DYi64Z
wYQQ8R2xTONT8IyryBjj6ozhh33cFOAC7q6HSMVdOx+538q2M2CY3UG5702PnCjvGdclFiOZyTnT
lTRMsaRgsnur7wSHcRGfP2BoxHA2M1Q1CIw2vZFkh3yOS6wIsN3xDgb7LNVmEK534Rb7RATrjpm6
ekoZrCMkbb4QbCVl34u0SaRPoM8yiaANkFuDS0DmUK9Kn4E+j4FzBcEDDi8HjV8gBLrfLUDBpiTb
/gv5hR/oA+p0V8Ty+4OiCUk1d7TB2EJo40+hfK/B5kXZit2okapfL8lohg8gzgt8nz6R8fVNbzH2
1DMwlpai1s8TJXQSLUDpMAFS7a3NTi35fyFDdkaHUNC/5k7xsYva400PpaVHNVOCHRf2Wn4+F4Za
4BLGGA+HSg4XHKzKBKZG073RocJ0I2rntooYiiN9F3pZ84hH/6jyrf4LP1jkfMF0PrTay+OCgT2z
Epjh7yZKg/JaiZJejpvt4uQqzl05mWoeGmJvTNlYUJHHNC58mw/C7bRXvry5RNbk9quoc0KPgbRh
2DUHS7KBdiOMBMx+OgcNe5sE0f5UKj36d2gM0R4gLpVuufIMtZn+CS4nhotw7Cdis+ajwZdDbf7+
jgwp3i/WE9WvPH9N/PVjyw1aULMlmA2pziY8xZSveE7KsgxUXxwzSYfNxMntolmUvPhv1kHTF8jk
ZtAwBUiQ1LHgD10u1aCsCOk4e6mKHMUUqrGPuHZoJ9v+4d6uBMcN/KldwnVN+eU7AXSL65CCB+mY
LMgF04tX7XTHwPLiYqUDHPtg3qtRrCgzLD8QGbns7ozN1Tjhad+lyvwO6OpNG1M8fBTF3R6MtvU/
dZTXwl/vOH20VqGC/bhGZg4g/Y8eFF841mz47DTTjrQ5gofK+uPbzYI03zChmc12KN+XNt9g7rJ0
OhcmEMDR740VjWD9IyC9/HH1bS7Nx7fqHGWL/xV4lECR0uF5gCETQJsT40rlpmntx7Ev2Hu5lORQ
j/XzEcqhGxxeOZ/NJb2jU/tv7rvZPdy8/v7r8zUsxpUhOR2j5ckrx8zaS43wCBIjZl4c/NWL9Z05
epVirJWH3TXxAphTx9fw/JUYy4XjpQ5MV/DgSUOSaHA7A4avftvMWQNBCtxYZGw+KgdvLowgWdqf
K4XlvTMQUKvzWggMSfAIiZ+AZb1R6922EO8mWuRPYN6k1msTlD7JypXfrF7J2tyCR8NOniiqf4Qz
t5rfZwG6TYG4pnASdGbOI1hsC6ucK8W2xWg8zQkkENTS4l2/y3NING9Jdw6hMRf56G12gQvJGEOX
yvWb+EWPh9WCZSYwIRyFChrgfbXd8njPScdZdWBcOumbwGOnVdctaflOrDi5kIQ3XfrKJ+ATdI6F
4ix3ZvQ9jpUghI9bo2iijec1kVgVuVCXW62Iagr6hiNeUSUh4h4kIxlX6RtkWt52YIZAFYTV6VQ/
+QB951icaarHB2MeGgJxRRH4rXTRe/GIIRxvb4V0b8ndlIygGavOHkXfPYKwrawdwvBSayr+BJqf
Fr1uxhvNgliFF/ZkQF3aku3vW6F1w8IIO/SOdlAFRRfGWRbItBN4Q+4t0htuGQ6FzMJdTlDcx1A7
P3EKxjmjos9zACfsvsdKOR/8xXKAgBcWmrV07tcYUpHxE0g2GDqOMV7tl69iXJ7RVoy/QNZnIqYx
k7lYW/8Mv/lKrYDCYtGe+yM0/O6vaQUNARvluIhmAB01j2bzLuyK+324zEwENnzW9/4yP3iEvWNI
Hdr3XF7h24GBXsaSB2MNNKnwb1yK9+cAg0eLuR9qiCseo58fTd3uwJ20aVw8ZV0CJPKJECjYwcPB
DMhWCY71LYodGEazGqxkLLbjFPg+1MiUuJ/2wQamcuqyS0pXs3QwHudk6Lqq6Vr5hKInDAenjwKe
VAcf/CVhqG52pHBpGF75X6NG8M9aw8rgv/VGOiIAUMNZYFFT0cbiFqGAm1GGsa1O7Foic+/XMVXv
RCvYz88QEmh2h2wjUV91dXoX3w++/6xio/s+peLT3IrPFBPwyhk1H+GQiM84IBrUoGZbWqq1PC86
Uu9VXYIXa6MYyMrXoZ3UUH1ntXPWgxxzloGY7d09R5n8tiY/9iLzGrul0w7QJFc4dQmYrlRL3W4X
diNWQVB1K9n372E0J1h1mn/tt26iQZXmiyfaf9Im+P4mCaWR3zvvkJXcP2lkI1he2YenfXMsUDf7
d3HhWxkm/1FSA6aMYbECT8EFEVCdwcyJaPCfBLciAFerzPkIoni8ZjgcwhzE1kGarKOoiSIg9ybR
iQsicny6A0MlTMIFLSlBDh96jIWgdWG+yR3f3gdP7RmNqtTAwAIz4oi0yEPTiTVrmPcKb8b7rwjW
waP2AaBg2Kva7MtiwQ/1hoEVklQ7OGBApGPz+AWfmdRZ0PcAt+MfvsHx+YnyAwvINmUvwItJ5SeJ
Gcx/sXGhoN8xL+poxbniBGXtvSDOc0t98OfQJkP1ZWDgwA+p2soI7X3w6Uu72CXLjqDm5ZL9vT2O
rJeLHVXBvoVoV5VsKOC6r3ZamQBIpJ/xzeDAEDn9dfilplRuOgoB22wjAnSq2BOUmZaxaplbajMn
c8sbV94UEWIhJPlKREEfVpfrBzy5djGw16OvZT1VNmRGhp/a4mKpoexuFXlOSdAXFkFgdWlRyF4M
iChgL0Jn4ECQxqOnus1o4hfC27kKYHO3bGnW9fsG2Y/stxgcZqc/JY7oFuocolS0y4MJD7U8S0X6
ZXlbK/3smjN0DWXyz2353mFeAA/7LidgsvdkzPB8DA4CuDdV0vJAu2PWJ2vEadt7iN0KyQcQaFPI
4DuC9v0RrNZILNV5jzK94/JQt+jTRDWsHSwv6v/hFIOZvsbjZs1z4lUxg79z+7/niP/bXjd1Ook8
dVuzWS2MCoqxZwUZMWxNTO6xkLQhxC7BP2Ku3uMY1Ib47apgZsAgBvkj0PvYdQtpfk8+vwMPL+No
sa7cso3bFtHcdL9BVZ5OY1az85vnTdEA7U9oh++cK8cPDWyiuLJcLcoywdeRNYwjsYaWwTJlNdMU
OHZc6UEyohJwwbmQfpn6BnVzU7hS8FYeQcwkY6osjq2FhRVEH7OmIhkUpuADsNfH9r7WZaXReDAS
rqxDjzZbfFx4N/qnjh/tn1+tyGNN4jRmwoEqIEdEGzBXwC+f+U3YAs/DrRpmLv/8WQCblBDVgKNr
LPx3M07DYTzWyTtjsBYSnyNALqcvwJWmxzCD8gJ55yaRQEjZuB8hEGDikJnTYjpe8FFp0Sm8ATAQ
+Ag4V6TkBEaqjhIIxTeEE849ftQYnJa56M9Eeb22U7+SPt9YNYJD3Tp/EEO8/ofg3bVBTgPVfAlh
n3eoP3hmb+WzmIETA9ezQRw5/i9dJ+owhwuT8tVjMJpmTP726yOmfwDV/5+phwsQauA8nj7V71Yu
Vnk/5QcMXh3slpllCfKUqGPXGp/o1QpbxEd+CW9f/jrsMOtRZtJQnxaJef9x8xMiI77zN1bhO8LE
u9IXtM1ib2tljTFBD2Kjy/Bf3pt3ESjaIY0MU4U0YJOLJxiqRZitjqduoH2r49gd27XOmC+prwBt
8HbD8AbP/2qbeAmN1AITITEecKwrkrzekSfo1VxNNcETGLp1o7dIEnnBZhkoqoL30aH0PJIQJCL+
aQ69LHKphRyd2yV7cLWhsCAzP4dLqjfcimZdQQGT9lHDAhzpC9qME1/zpoAHDffUf0m4jnjHbsPU
+k2zRDEB7QvzOOlICWBkAwBLvNN9u9N9EOCEX7ob6B+cRMw06kkCoz+3wm/LZcwzszlEYG5qGyEH
8zGL9m5HP065M2x2MR/hrrfzBsiRB9URyrJGo3f05drj2bP5AJtjxzipWfD+zqGMDe87fwz1Uabk
RcWZiU1lQ9lA8yDx4zSZteY/mCISFv+X51GuwzJFJah8NTfD+3tYaizpggG+wlCd58P9hAt8m8j3
i9QyHX/C9i+FS+4Y4Fin4tOCvfh77i8N8wNTj2HAWmuY4gLf10Ii7283BtARdkEcCKRJdwnyWI0b
ot1i/zGt+OseCG5skk4nkIceM+LHrX/v9sR/h9az8ZeDAWOcK/lgC8DDyjkl84xt39Pkc55OqKrB
XuhmidUDpyMEhR6MuomlvPlW9h44/XjbzsVG+ZR04p/VQg1Ka0BMVmRWSNd7BxlphbpCo2sWEloU
M0md4ysUsObEDhX/ccqPa3FEBgH93R7RwwNqP23Z+cxxuLr/aQ/ngV+Y9x/Rvn+s1dLo8q42/NGY
+gJThfF/Kmw0v3PHwuog913wFWtTlKj8pa4zeyrmdVz/a6IHgunJyFo/u9WdeVrgFkv58a8aQxhN
8JCkjc5KfjWx97O9YySsHF3HQdrgzqnlaCgv14tTG2p0ESMOnLmcHCpJVyi6zmHNvvAxvzSSVH3E
7n/NAjVjwB6BHbPcPxo9tyJkNveiPtqZ+1imlFInyhNdqeLFJJAKLtx/q3MueyfUyIW4H00qDrhD
wm7UknxDbBke+jjK30BYMlKmtsUU2hQo2TLwv+kGG1ChWOjukz4BCaiVXEHPP8UIeZEJCF8kIvlY
Vf5BgFUzcGJj23t7fAPdsEbg6iQJgSY6zmpunhougHDms4QYeNFU8lgJE2+rWxuhS8GT+E4yzsFp
ajtFUX2TexyZVGhNZedErGq7ajguw/kc1yLzWPSRkLze341uRmP21QsJbmYwb3LyP99m8e2zffZd
nEHtlRl7ua9DyTudmcUqlZKBgGNxVpY1jNCls8m014IHCIPEtAdGz9gcG1fDqAlSJPl/ZPfXklKn
kz8i7dYCf/2PKuzTiZv7fjJrADttSCaBitSfsYl3mQd00/Yw/XPZkoBRjiG2rBL28a5404QYGZOg
fQQaRrqi00Kvp++Jo688qipT5xRvl/0JNP2gxlK9vv2n7mGLA/WcqGKofHxuubJPfkA+PJjd1O50
yAAbRvK4frHn30tT5V8UBk97msBsQ0SFE5SBnV30i0SXQga27n4NKkoyMWx8ruaLp7g0gFbP6wlk
w/AjEzQz3XaEu42J2PDH9WDGEAzIRW4YrghwtjAIm4BNgyEtN/Sgw4aDuQ+aFR8mIVmv00qKM68k
l2C4Q2ZHN562K/bHDNYkKChV/2PT5hR4Vn3wn3EgZVtay9Ykm3WgMcM9BRr9mLTkJgCdGThPxcUm
I+UACWuA2j82L5W3GdLDxURJAugXHK3IGI+m38J5CWycEsJGRJnDtO3oqZq+z1K+kvSHUqwrKjbP
O7gWBdqHd0tLD199/Hj+L6yIuDI4/VBdY2rkDmwf0M9GCX3ORUNUk9YG4RvHIWwCZVrtl4Gy7Qqf
dEklgb8IiDEHSUKbSQPDhD10ah2ci1jd5HDH2rkA+aGvrLptgcM/PBZTvR3k0scN9Au/BPBH8kbA
5Y7u54N/s5zBX6hDvocWU9L4zPy5h9na/ihHtMXiBiP3ztcTwmd1VNq7AbnDKBcXQngJoniR12mP
jr/slrQbdwIRgbZ+chWzZn8au+BxYqD9eMnqaobOup3hr1AFNrPyq2u3vUjOwiCPZ0bvID7CXhQ5
jhrb6NQAeGbOf3HIC9i9Rt+XAxcnosre/xJdKI+bDoZ9Xyo+9NKIP6Gm/HuAeYcZYODfGAIOMBjP
gaaqQyfxTJV/O6HpRT5oTr3Wnz19ZV+s6L6xx91XC2MaleOYVFXDen+hbXb0oU4RM03+vZg/Uc60
sdnYn1ifR/yRACrKDbFmEusKgv6gYfbiU+g4Lph4LJ2SNOsmW/e3C97eB9sz1CX8zrGkgmGiwWJb
q6gkONo0/SwW9Mdp/OFUitr3vZ2/v8LqpEJ6oK6a9vU7eMX9Up7nPCOXmxOUtji2gMX85IVGrmrK
OkINtDK0rHdZBG4yoLm73tUb4ODhPYCRiyavqAxBg+QuHB/iBhwBN2QZyNWSRJnJ3av4yNqRGCIo
BvgWHN6rev+UW36IzA5G1FGbmmGWi11rmfjTjNnLelck++R3aCyBACESNXUWPytHXV1hqiq2tG2u
Y285RbeQwe79BrMWX4iU3wjej7InLnEGEWgZphKbMvmoXlCPHqM/ay4ivpn+mi6SibJHHqg9CzYA
qunQRf9+4zVfIA8GHzt8a4Q/f0HkDVvo2oKTGOO0pgv/fQYhTmtSiUWua9Rp8ltjgUm/NIWO93bK
9e82Xni8ehO+UsTciU39wqmSJelUI9aD3P0N6nBa1BH/g0x5mubYpBHWiXKuop1g30B0DOMGrsmZ
KFefYeExxmkiUqRf7XtTB1RIKYWDz1wO33hA37s+/Aa0S4Xt9JWrv2fO/PZ31Npvz31cPyDIgq0a
s3A+yqXlYBMngY4ZV+vza7SWxfkFqIdDnWvq0mjKvwQ/Y4DGbZirtLZxu80WXlFOblhPvFW0d06r
ZKJBbZqoBa77blEaSVR46q4an1io3sugfH+32x2iqY87m3uRMTxHFJ+WgO/rE/1zj1fwfSnaBYvP
kbe0bDQI3n2wcfDIOw0tZyhxH9LRJeOw9yHjtZpFO9ZY6MCvWzOZrjX2apqqff+4Imz65b6+XfDr
hxhL3HZVBVUvblcu4vk0v+sYqPJKRULNDBBOmMZhEuc3/be5ltwSFz1EicxnGd4fjyc1/VGwkEDb
ohzHRTdGtNnwJce2Ml+nlxU05aLh1U007YJDVwcC5aQTvXYClJ47hhM1raPMYbiCNroKWgUIyiMC
ayaSHOd0RpMgHcWFM0VxgGGtbn6X1DoWCHxHhRNxNOQI/YC1YizlovjmxSB9T6Icd9cor1wUmCfc
k3kCIYWwpsi9i9v8nKuDJMZ6Dh9MtCie47oCfD825yRW3IN4L8Yc0WEKJXtJOpwlT61MypRaDtHE
EI5XNp6C7KvWOl8ahwz6/KIkWjpumJMxTLvSU0aBHirEj3rTE6/hJtSTC33u28Z3tEKRCLXISDQd
bkPiom3QLkitJnoS1CKE5siBFqGxe33VFltAdgqlEZiaoeAOKsBIjrWV7jb/gFhSY9dahJvebN2Z
IhxViYqlzJyEclYVEihRK60lqqkXl3OVK/sypyq17tdhfW4XAyih866DEgqi5QXEoFrCCkhKx4w4
IqZQiGNWPZ8HUK0G8r5z74fdQc3QaaXicENvv4H5RqrrIuYbx/TG/z0Ets3Lpl/rhywEdHLdMkNX
kGZO4vLTHLpMvsWluusTtXekR7jVYH0jhTvc1g3NhfBLabRS+a2PUzQDLpKyyxPtaPRgtBqmOOB8
R5Lg8sbWhuosCDb4KcjNQnMuNVYrQoxtoUrzq7KpkAMCX+Tzc8Mqbe/iJGpQhvfDqZWkezWQfLij
i3mLK/HWkivkCEgUEqxxDruChodksvHQJAsn++gPvw2uHIGscijX3JAZO5FPRk2gMPEkVKiQAlHA
dC1CWzE9gsv48c1nnJeON11b0r+nCPARtk0aLmS5gGnhhhyDvBgApIT/UR1AtQM52Oy/utZ7U0nz
MZhSV2SMSxZNXltVqdrTy1oIUEDsPzpZ7Qi5eL0tEEGSusKhD7JaZiMNpfPCeNjfy7zLwBW2Jv/R
u+rCz/s/7+7zGrNnWZaQQNtz5FAODav3MYWyNgrCowKSxUKsbYIqlhc3XDAeraEhHc0FKuHtEyET
MgnrGswlol+at1AcaFEYlbaUiK0cy73f11IjdjYzQt3qFavGt6shiw3/PbApSLFsWvXtz852Z1vk
rPs1tJbXVqvIwpeNK558vW8YfNa1OOmF/6lwsPZ2iLGvS+ekQrU5GyDZW51JmZqDBfjwdUQze2sN
kf4VuhpEZI7UhGz4ubr1GvG7GdVO/ppwJCtMwzZg/qDNxK3u/CoPxgr+kJr+rtWtrAkDoLw8UXhl
umTYIQtlGvjst+PJnZPxkD6r9FFjFlfSqLpTN7uU7h1dxgcQxCnd7s5MUriZExpJwVTXZIBIXTpW
Sdi6D8eZjD6J/OX628MsdZ0Tx8lOUSH5qp+G19MHiITpZn3lyPu0RVesAU3eMXKJxnC2WzHZ2SAv
/407h+dwTdYdC8Hfz5v+BPynwixhIGr8IibiqsOlHUFji7rkiraQrD9GfFSTadwdV4ipVNiBo6ca
vV631b+NZjW9P+smqwgKRneP7CHgzZ6X4Jf1GwvoMjECnPSPYt9sc13hzIT7JVUkJ99PCHtv2LPi
r9rT6Fibri2z0D2F2R5qx4lICBVUbiENzz93TL/NKJyWNITWyZOp2XRPfVk5nMVQoL5xkz4HV3tN
xVs3MM4AvXNrW+7elIWpyXNcvBu6oxenogkEiCAxFOzK3Sa1XXlQWaKaS3jrpyeVvZddH1uiDxj4
ZsXRH/PrPWQYO6phDLtHuTOWGRGoD4H56N5C/YdLbJtrJIBN1nqwIE2rjCNS7fSQkdIXeVI8bBnl
Hu8JD0aLFEEJ2JCpRV2hrGkzjUwDRKqV2zr9/MSz1XgPje2QgHugRwfnFY1+O9xn5aizLa4xTVrN
YL4RAGBdzgk3BdlMVDruXzoxb5yD+FEQz4CR7Zi8gAKgOeGcbCAYfrcQiRwaL6Bv/C4TQ8NUVE3M
LO7MdUQ2diRMlWm3PNPTJvR0GhSUBWQwPbyqbPbI9yW7QMnnOoNWrdrBV6bPVIOOqT32iKseC/v1
+uFkJQDinN1jz5e0DxMhb+3FwXW80jpaSkSRc/71VXHlWFLDHlWYmg7qEoVOtB/cwRrXjk5uIfmB
+S6zjbc6CeZqpScXkQQ3GnwHLDkfOQ5z2ie/4Cn07S6ugVeeqatpsV3fIixRYCiJrFQAtKrQgN1l
8qoTYDqBuFQ7oAMdHHKS8qa8H8cWtVSEE8DfiljwZeZtCMAfOmjzQ1PIq+m0fL8P+SmeJ9nI4b8G
4EJSrfHcAu3Xk64gemNo+nqErKWKTmyxi22z6dCyJLqKBi+0hqiP8AgXLR766M3drBcR4S4/Tl8T
UDHD02ODIFsezDWZbdv1jw1LHDMGpc2p+UBiA4sdSs8surgx7va/meWlefJHDmVFVE4Pygau7oJl
ezwbEQkcsv/CddgfjXRawMmhRUDEcEs03MLm1jWk910OEdwu9aFTCgBWaTgE+Cll7xaoiYroYLcv
WFnOIh42TOfMOCSXwGyQg21iQunHAyG8+TTksCV/5yK4tShfGOOlvgn6/FpukZU4X0jYm2LPu7t2
b7jVplVfGXtaUnBogL1KVyd+ViQBn/o6nwazoqm0CK4ZFCxbuZokUdTTO7yNtszMMwkij353QGFP
HuicM9vCPLWf7m2Nmcf1SBk671TTkWw5qtv3lufyHSVjj8j8KrQOMHZGSe7XNFSNhTnhoteofu2R
tDYuGIck8VnHFpLj7tYVWY1RwPJqpmnzY1aGTRm/fD3jZL1SoU+qkIcedD/3fX/XJR3dCdHkUD8N
1KYIs/3hz988KqMubanwwiLYu4BzkMqkXSHTx3Eq41SLQSXMMxuvRotnTtQYKOne5vi9GncllxaY
HmEIP9yfH2boT3D+VO9y4wuSDV1f4B00sIAsm6lcJ3LJ/2Zy5iZvyT9NrkL5pz6IdBq19VYbKNh0
TN4t0IraLNzeZOZxY9qhV/7dHdcBKc/3sfXBxhXt3J94H/UkBmKV2I6y6b8sMUEbIexH4X4wDyJE
i/Sv2ic+SX4lkMwRs9ISH3QQij855lJRqWN4OW3nN+r08OfhcX7Noujt539QSQTPUYmGOZ1dszOC
i4jajCZyZ5A7QPGkvVUl7K3dwhVm05G9dlIUWpQzUM9FHOVPVNMxJjXCJWitiY4Ub2pE3FDB2d5z
tRDnjuXF/G0k2nhXUsoM8lIY4Y0Sku6xBve70fxOWjmLEEWDyTzvXzUGoaZpIT7ohtifR7Pp4MOn
PmkE8hTHEBeV5CE9QUD1+2Wve+tK+UsKX2KolO8O41wWnnkTeKBzO6QRnd+wt4nOFIxKqhSxDQ/P
QZ6N2ZPHsF2iC6q3sBUCtKufE0GW+tjEabjF7PoQrviY+D0CeP1z2E019NXofezn1xP7423OLyau
CNHN4pZyLNt+bs2nDWndEYv+5571UAtqILu41uIPv4bhv6+ZfS3x4QzxOjRPid1WNiRW/0b0IcUl
B/Bdhz5rTL76vfJYyjUcXnpf174gduzWiQTkkvOES/ei+Z+hBkK75N5V1dx34hKO1pNJSxwT0MKG
L6APZ2ZcA2M9kVJ+s0nASRC5cTwwk/A1f2/yxUqQSJ7eF/fHQmaspVQ2BdF+sY7Fv5UdrWx0jT/5
HA4hmJ30UBHcdbef3/k/on0R0sjqg8hWPDdZTjOQ+Aoc/6Srml/Q+t0/5TW0ioFxiIe4O2L9TSXZ
JDIBOlDXdquLAzwYPhmPqz9j7YjHeiWe49q2wOpT+EshVSoAT0voaHvfM4vlgBIxEBYuPDf3Elw5
nRkMrE3PBF3+Q11vZx7MaSIG2MH9mQT3cCOvlzrxe+qSuwcW3Hn+93gCB1EeqAzh31m/a1sKHXb6
OhqPq2K6xnvZKyZYxZwtfA07LHbe/SauqJ+Cft/OtSjmVCvFqplRfx91eRDVflN3QoyoKh+WF99e
Q1H0FDIdDOszDsLU1YEn1ML5E6x+DFq1T/6bBWkfsdg57cLuarpPz4toX9s9fFV2u7zooIl3GnyC
W1bJYqqz/71NyWVPDjV8FLLCNaYJitaK8/+c7Ja79PdzBxOZGwl25vlfOsU0fL8PTimW3/JUP7cv
RtDbc0zBCVHx80xCYt+AT1p4hgltXFfH6qwzjseCZEqFhKjFPSDT5IFycC9UiyWhIBiC7ZR8nSmb
LVEyolL2jBHWylVbsyKMIDzvn6BD0gPSa1+4KcexGzxfc23BoQbMwqDyC/R2mCwX+cpcKYewjBnw
hKcfUNpt+R3FJCxJKoeVtXifen5QR9cd2oruaY280JrqPVhc5klOO1CDZ2B/hT2JbGSBVSDUmIxY
mgix7YUUifPRx0Xj41t3/1eUNnjuaNADE/9vMA/dlJpJ4m08N/jBqjkiCW6++sxgRdw837JwopTi
ht03daMa+gDOaQA/MWMqZaVs6yBSITL9v+VYeHLKm3BSVnnQSxYTzFVSO59p6v14AV/41LGkMAmR
CTfg5IvtAJlQ5ZiMJGR1Alr9ay0OAcowrv1EtFxwYlnBSo8hL/YIRPDtA3/FXvveBmOG6PaFayQH
HFEqTrmCCpYVfKTRKXaXvldGtMPcnJ+8qAqISp4Wc3TO3mGUha07WFMOL5+OQdgMfU7+GMBIReCH
lgaRrexDxIBh/ipiBjdA9Y5MGim2g1nAZtfjiLqsfhwxt9NfntakIx6la/h+W11q+9nBQ7mkwMtQ
YJeC2n0DshpqhvqE27/p80BcOj8UV2oUHJswnKEUQGnnLe4mRndijFzVgDULWuOnxquq7bAfc0BG
aDXwbhP3w0IRGMJ5rOWiq49pmXBLF+A6nvngO3hLDV3aDsmoAtP2AtxC3qpz5t9Do64ub5C93kmd
qZUA9cByJR9EpAKARn1y5AOD9We174GDDIKk/NHA6wRRF+YyvzF6QoIDZChNb/kKxWwpVij+qlWg
rz7O2uFIJ6zgpuz8w6gRZfPzHvIHVeejtOA1QL439QvX70pq78D7/NliHV/jPlgvTUdW6DMSvF1R
JmnY6Xw/3SLH75vGa2PxiNCO96sa9Xu+nY9GpnMVCuveZIYPo0UDYrhY3mVdgQ8kpTtLq3nZHTAx
QJ8M5zjPz8nzrdI7cojzBD9SKzlTyDC37FSKnjQeEYcr1b/KEa/CBi06MRdhpsj7mDYHKKQFO5md
G1ZQ6g01qOkWwYGd7uw5CfvlljsjhG8rctHK8bU/fN9pIZMr3kdFpGZgb1LwXPAN3U5j38QhtI0Q
ZDSswCY5p77def4glfEoW6MSL2qsPTT9Kz5urh5bbnLCmtpR4ZrjfUG8f8e1/VW2AuMy3Xn1IwtJ
XszSxIr9S4DJB1CQXBHGs08PW192bbHn8MTFRjfm4uW4InK9XxrlRFDrFLjiFFia0IFwGYdB2V7M
22sIb3E0l6qPhHklaw7eH5GSw8Z2VXxUaHjH9dKFsnD6dUbhcx9UuOt52c4eo3uN9eFei133afFI
K6f+TpihDwAjeWyR020O63FdcJ8hcjVxyLBK+Qy131u89SWyiPwJ37omhMYtaXhMM6SoSlAKueSL
hPawLD0msS31ov6nKjKlrS3LfbiHPSpPS6iocNXX6dnMAZUCtnabf78gkAByMjZkq/JNtsgqPEQv
zVdZKAtCPujII1od/YOstpxhxy+gJaG8RiW1UZ667n448Xo3vFC/NkdUN9ZzZwlSQRhimI1IwfdB
Yg++YZRZImKZQzR5GqEI3G23ptZsN6kmmJe2PyFApEzwz5bUV0FqpvI7YKxlY1ynvWU0f3suXf0u
02L8bgmWB47DN3pM2aMQUDZUERW0VE6YurUJMZUPq8k+bh8pukPiLmHDBnOC5nhU9XktYX8zNh/E
tFgvs4UE3GWVz3k+lvjgTKeccFnpyOjNDdBW/F+ytuAclKcrvKTpn/kvRakrcwxAJSGUWeJjZ7oU
XL7JXEHAhXHRjHbBGJMAqn9MuOd/9DWd0sOcPJFOLE8+wiA8sEy7rWLn06VpeR0oBvXCbZggOtNK
j6bYfydrKLwU3At8YGjPWJetF8QRwdFMFAqNty1PYSC5CEpwzn5ysmAG3n/yLjqBhovUrLsVl0kF
hAg/wGpguGrUb4K8UByWNI4qVOz3liiuTQWJswEFUR8+etvt/HwkbxsM/a3/X4sKSHyg7pIDAf9b
PSqX7AtXa28qUT9r6pQSdTaDhgI1tplRDPbt1w7omI8kRkHTtcYukq1BNeZKOBoUjpVQN/otRc6I
cUUyDU5sw3K+I8/XBnyvHmWfQWjc1HHDyNQJG6tM86FKkVP4qFXrzI/jipqvHPLJTU2p8IHxsna4
EEEe8QS6/+38xwT22EmrHNBxnbQJR2VPWFCkDrl3eGE6m2yuphjPWMkE2SyhpxGjE4CLXqXAnifI
/CS6mpAaWjzGq6WJP2BXhzOCIv7HRKCmfkft+C0t/sH4tqEcQvmi/snQsCqXAyV8MaMrnXOcJ9DH
sGywc3Fg50ySZ7i2ZTVtsO5VSIYBtPhqZWdDcs7xxdkNR8QY7xlL6MGvfggZHP84QeH1YecbN+h9
NgDuxW27Z8dkTQiFOcC9ITN8LrnPuDIySTU+/TaF9585d0V+IBKgQyiQmxnemyNwzMH3O88zbfbW
FyX8tieWCMtDGJzfpkImdb0mtZb1iaEEZ1G+w9YWJFihHRv46ijJhHdYcDxeq3NeP1Lb7pWiMFBz
MVG7oarJ6YjccPC3W8FlEAxpVYmkocSW3Y3fbWgRtXQkbvLyrHzHcQI9r+ZooPnfzMEhYyqHT/uw
CUhdXkt4UAMPRw0QVEfSHb2WxUWVcDt+x3V2DLOp+CStOKHL5PtEauDqZXn8lfkpB0kMBv9FTXYr
U+gwJ72zynIcdPcajDxcYBmIZCjPRSQYcz5gaE2Cnlm9WYkQBRX7S9nQdjLailY3M+culp5sGgJR
bT0n5p9sS2KHqFg+JfJEdeUqVbldkCRlVOCRhksV4PYbPpJnRXMq8DzzoLCuwExIUleFl+7UMOp1
On80A9akrn7mO51XlS9w5HifPlKi5wotaFBNYtqPhkj+AF+eoqjqyInA4rI3tbbM7ALG8k9bq/+8
7HRrZ3WwIgPH4GxNBV0HRiGrZcfdsTLWFluySQ3uwP9GM6MsoKlc6OWefqQUjWjXnLFb4JBSch6+
GR9SVo0lQd8BlC2tw59Bwkc/eczQLTMJy2015sqOwe5mQsPuXjCvwdS8S4YCostdUgf2kJYgdA/U
8yh9thv7Xqtudn88YNZmdpi3vTRo6DYSG9OumW7mx7HRUlLg90m7MXqWF8Qt8oBYTlomEuVj3gzr
TfIDVQrhLeNutGVRPRUhHxX4UGnGBGKwMHjkgJ59t9TeZUVRqcv+gwv4HZYyny4dcHfI/ghctEHB
MBLfYrB2M7a3oIGdjicej/0FNSRmFJwg2ICdGiKIyWtzS1LEa9U1Di2NI1TFm12vvKouxAvUG9w/
QD83HAmrDCZQOmM/X2aAm84WcFXqYK18qGJdqgaGqzhkgAcU307zUN5C419IYQ1zlRw/zcklMWFK
4ljR6LRDNw6v4h9FLy4PYrpWdy0JpgKGfEHxhUArGiovpLb4T/ryuYG6yLx9pUf6YsZFa24cXrvW
6zRzJayl+83u8v13tCHVKjdyn5VMDMGHGS5ULFrdxahAoSFk31OigsuL0cc6dulaWbBI8yvYa4nw
FUyxmooYltoy7O+atmoAzO9TyvVmji0UOfRh4wiD+v6aXEplMOKFkn49yWa20RKH6NvR4///VEwU
RMI0DcxE2eYvFeiROUWuGQ6xXipdjnpAUnq3G41m88rQjlhe8+GvmvnDMo179sh1nRYVv1/zq9Su
6lJRunCG+4bEahIAj3XEKHWsWgHAadj6Z0CVIG6oiIUFrFI7aUImyA6q+TRgLZAvWEpqeSPEM4Iw
eE9zLkKJPaA33RkLMR1KiUe8fN0ECgkl1MZ16NQ0mH9B1uXPFFtlNF2QN4aWjhh3rnfG8vB9mNEH
9hMU8AD/ZIYknle6tBWQkAxsc2rPNMglG27XNR47QaIpX0xhd4zNgc8DoGLILEgIt1N4UX/8ngT9
Mu0MzZ4NE+H9m+7ET4DypI7a2aZlq/BBLRvasnLciHT54cMCr8I4dd0xmV0fhxK007TNU7TIyLhY
FkM0YVixAJBwvYyWdj56H4fJUL4sb3qhrxUucsGD4k9KKDpHQCCnmtwgXNurEaPZt5vPg/SkKr/p
vETZDFbyTgMWdB5GYHD8nCL6aoWqmaT4mVMD6j/bhUxRU2UJVoZ6PQxHT9J4mAH7I+pArdU2jQBC
w5lcUPM2tEtFrlNYIjRhLRtyR0ljp1uUpd5KzjVYGG3vSjwrrItfiBCTxCa6LlpxZsP7cMTKHNfH
i6tf53c3WtEkxalBtH7LNcWVh+bd+TzqafNkU6OCUTkexnLgnW35/pduJ5J3c8U3drRT9l89By0Z
l+iwD/CxMlnxtyyNCj7Lpiiip2g7OfTGvHPri+gu/utn675DsUNRLEhEkuaDcjCygR3HF1HuHzuu
c+ryMj5Xp7RAspNdOEi8QPePTcw1hHWyiC2YxCRra4uCAWITHd9pvGqlAav+wWMv5seStQLaPH0c
Ht5JX8NyVmrcjmab8xc0G4rGwzqmwDxvAqgulvcvuNQcp9uOhul6CkqSdgdRVf/C8VIh+47GbHpg
GZl3hKTQWvedyg6xp736UjILn7eD/CvVEAyeNA0s/rWtHFRz+bsD6ZRBy+jOavolglxyuOMG6x0b
FllYWkjVckB3rKOpT4CaUyxnr4WfZLr7BjF6GXxEySeeGHjRVzinaGehLqg9ZHe/dlVRbq17Q8ee
+9+YMIJQ25S7JjjzALWUQ840Zr68A28/sEB5r60NW1oPw8HtDLhq/EJhoMrwanB3mopa72EpVeOi
SonGXMkcBVIhRBr7kp6ZZG0IioDIQFIbHSlPisQn5fDhEsjFXqfrRrW0DjjCAJY4XZDXxIgTEVnK
WnVBb789xlphKAjFQgWDSxUz5pr+j0N5GJOKUksJrMFSyKmBZjsDMQyDoY2O25kpv4K6Tq9+2w6j
ZGOmJzZYGAvcbHgRQSUrOwoxVqeIRXczUyyqmIEhkCrJFOJFBvu+PDDTrvn+7XH/UexNMvhze7UQ
dn70KHix+OkLCq/y59Z+4mSJPak2+33G3hY7oKUvJHPVsnc2bxRY/er/wnuSKRBp2J5kvjlrZDAz
fWbuwK1NseN+kQ4qPtpk+A+9VDbPRe7vNLDFEV6CfIHtMfRt8jzZPqiGuRoCoIBT0XT59Ghrxs3P
jZwaFv+F0Tu1SmzaeCneoEByjR4jLS2LNZYpishJwEdVvT8C4yb7w2TrqQon3Oo811pkcf1/CMQO
FaigTRDoQX6tcaNcLlXiSv98DBZPTtsKcEQ/iiAlkVS9XvNiL63DRwq7ZgfSPsbn4O7VQZsKzNop
PBiEkcCRA/iPymdxAATS458MKb750oso/3R76ZOcGG3geo+0D3RNVTLw1xLmuW2xk2Ge7ok8CDB+
mNLAmMihLn7h4pv+NwnAG0cLdtW8Fw2D8C37fSRGmrJRWHjC+pLE8/kA3qMiVPM3oY7auvYKou5A
gXwiPDJo5GCGXNSnonOHcCbGujFSYR4g9SOjKnVH0lk1/r51S9BYCO0QNJyl9D20XK9tZxUSrIyD
bGGIM/PS3OgG9EjKBA8xMu+vODFl6sspmjbFQON3LK2HANoY2k6cnn1ThSBFCW9ZXaT/r4N7A+7M
SPEFVsCewNvb9oDqhJZOigm8aMikYM0E/6HvDkMb9ivFuLZIDRdnkGS8eVg5KaovBdBDuVJSD+al
Cnu41HVwmoY2ZsFdef8Usr7XxNoE7AKTBEGo9tG2pj1rA2U3UJPK/bsA2O+vyUluoZwzNvu8c2E0
yPVerf6zeC+RXuRmgWghxrQDHfPOgbtDEDrds7l8tgC7/7awbCSW2brbgrx+6k2c2ZyKM+OdLNYZ
lF3f9lU1AOe7t9KOtm85iJf5FVw2mEpaLx/NiqVCmqbEobwrnHq7YH2yeSlkb+5fvpWj9G66/E3R
mAcx64bnshnhbsCBWUi3j3C5FMDs/03BiHFcSvjAFbXIIs9n8kd/uY8O+KiQyq22dZrkbu3f1gjb
+MhBKcdN7RBvdt1D6CsY5Nx95j6ExoTKNmAOFZMH2hkKYgrGhI4AM8qz1XxcuPBhbtd9eoqSpUtv
gwr0Y4g/NyZM8cYykw2v2I4iIvS0lR3qq8WNq8kPb9Yqm0ac7uAZ9bs/D2jFVPnvYflinRt4j7u0
Sbeef7UOeA80r0AMLl7VUnzn6h4FCX5EHAM0+hwv8L+cHjFR/6YCIkUYFHAzXZNOLsNnH+VsmLDw
LkVD9J6e0aHQXCPAqsr0YlehepBM42F31y5WZI+uJiOwOJUj8OeFaarg6Ju6ZoYNIH2+fqD1hoed
vud9jzEJ5cGDDkICgVDxRdZnJcpDsCWRooeVPpURdg/VCKAAD+gcsOq6V7IO4okBiCgFRMOS7KAI
u8SDOolEsaY3Y/udTfv4OszQ2Rqt0PrfQGMuyETKz1reEwwwDfg9rFYqIwbnyVz63qpDahGO+ytx
l3cOQKGlni1Ghxuc16+TSSL3uC/4jtPCoS4zpv9XEbSMpi+DMRZRnQaUeoPNCx0o0ky4i36FwjCd
OWfJZ8D1yCzuBfBFoSn7OiUhqxPNOr54yntLiqz76SKDp4CKZEISzNOnXKrYKpV5pUG5XY093W03
chamMHRSgu9QuXE40Ok+XT9/CJ16Gh5hVV2slCEiZmL7HdcyRyb1n+S+4T3RQCoCBikkncB00sEV
WxqrmwjoupHZR4KuIhXL9dka8mkMWjD8Jbcpk5xRQARb7Ek5O6vXucsiG8R9Vgr45/uglcLrpte+
HntE+4x1m667n4jmBWMRzOBULBeiEdfZaO2aU2K6OAHY29M5NaXadqgF+R1EAQf/BHgOpRxDZaVp
3VWwR0cgq7wSwN4NlZGuKvrBrKQ1e3OMlpUlL0uzmm2+UqRbUUlQIK+XXr8u+H/zfxN53IBTHsj3
zwyPvQ57zG+5uDjBBfjZR70fdwoVm4H9TCm17xltWVEIXWVNeV5XxyT27PfZrOazp7asqHIx2PwT
h26FJ6iONs2Ez5LBumr3P+YyCMVyazBpe0sZsWxfaIhwpnUeyOXtIF+1pz4WXDOauJMeBhgCZail
uBBoLppTQ1pJ/pNanrHb25fkphB59TycrSC0iINgs863+pYOZDSrePx2WmtuWemmg6uRq02e96Ri
x3C+yiDymQcUzspVd4trHTMfC576PISr3lVh9oEwdt8IUGTWEGVu+lNrq2LW84ThAHQYpuR52D6y
6PLI1ynlnV6wDjSBO4+2FzQTwgwh+iJaBC7467UIIpCp1bO/RSmAOTstPRQAQXLEg391EJUnVycr
/9rxD1Gd5BmP1fCBrAx6OXvs5L/DODhP72NlxjRCilI9FP7Cn9CBWr1vBFV1qbjKwpqP8LBbhdl1
XYkXnTITgJe/VxYTM1ifrHHnOZi3G1XFbCjpKh+sSbnEWUZyclZJKyC8OGCv+2SP8k4etotItT5V
1HVAAGKiSg2o8z9cS3QxCgkpyoCaogwUFNm9wTgi1av61+flORppBGiFVCqW3lnxzvlGC+z/TNVx
0FKiFgquneC707yrcRD7itL8jNTErDGT/IK40XZ0FDjhoaea+fdGt1Luc3DDfF7uc98JmtvqwGiV
9hcTTwajvdKDqgQ5QL2ePAg7oB6I5RYLavgBtPwS2zdkZQhQnd3NAcw2HXdM3u/3w9PiUxY6fEPL
As54je1NokujDagqn3ArX3Nlio67X/JpLpJS9+6i86F0rg61og+ssy+2412RmPj2wBbHjr+B+mUW
t8ZQXmR3VLgveeIkfh4Q/5GePcqA8cJohs+YqIryKdHQWK+hkNYZ60CGMDWotvyWTBDzimv24ENB
SsFQaEiK7ldJVbv05Cn5k18bpLisXKVnPRIB5zGHd0fzGS4qaxm1YgP6KSS84xE14P32e2ktxxFw
vEU5oAz/5ZzCrQ/09Ppn0/Laqt/NPJKvUiIuFmfe4MxoZ3iIp1fqow7FoDtLtZDxlDW8vw/a5aLg
ntqo0BKNfRn/wQDrGZuLjePLv6Yr2fQ38p5Ba9gu2P7TgkDWC6cArFuSPxE4jlnTZy1IySGwBKn3
vzdW55xE8CBROF0bq+ORovaB/SJrb7UDIlLtQv6fGCieh9V2uFzr6Q/OOC8vgP/IP3wAXsclLDqz
mh1/eJTLrsQH4fkicd5Q4G/mvN7NgSIhADeE+r61JbZJ6bVSZu2MnZ/dPjzc7zkfAYQS2ne2dCuZ
Pdm+WrwWWgnAYMWP4Y3eoOebZYL9WuIh30cv/0dlSZVn0y3RNZEFWdkQmRf3v7OzscRARUzln5aq
p/hrUqfTCfFrZm/hma5dZx45Ef5BJ81x+YJEZ24WsP3GbIKvzUcLw7fAqYp1KkaGmNuqssaU5ubn
Uqtrg07mfb4q/DSeIblQ8A3eYVBR6Cel99RdeCwQ+6hvrjlhPZyc6LdWfiDTfAPHGuGE/VlJCwKs
fC8Dr3DYcwEocTQ2DyYSAeva9TPFLLUvCJoGYykInYtWVLaW4VSPJCq2C0jKFWgHF2Nt9GeFGjZs
IKgdx6mbWeWhZ33DGNS6yf+4NVi3BwlJ5DXSCz4Y3HQnlZL0tF2340NaC3dzhZR4v/lx+NFIFckd
8XN7xZ1qydd8qJi7UQt3CvDvrIHOmDRAazEEa8UoVhKckr8v8vl/E3t4U06apiQW/mDlQkorli/m
EPgIKt6xULwUn/zhfVTyOuiojIPJ3qaoIu/za7U7+v+OUfHfvsHwm2Pp+e6AxfkUNLrqoHQXiaaf
nK5Z7DqyqFE2wlVfdmhUKeRaD4UFfFKaBmqlZd6fesGtQY/NZpEu6/9qEnRVqfiAIyaAIv98hQzm
I+/K+8TBFlUUXHA79CgqyUzTi88ObLKWbEs8j28flatDAeuVqPNXKlvB+vKUQRmejJc9afq7fptC
6lf7OavXPhgpj/jO9v4rghczhU2Z11gQHFFOxR42OSfGS7H2Z1pzbCCfhPBhbAGqXjk6SkPS6v+f
rcqIO3hyMl5LkuzWFFyQM1zdzl+zqHjKy8r+gAJU4M6ARkKezKNAk2qjbPB9cmVR+pmmZP/82QJv
x7J5rnO5dObQuYnODsbnZ6Rcn8UnV41RvUc987YgEBoRcYUtfziuyvLLdCfnU47HqZcZCrHBRrcS
nw6ftDxL0/0/y9GssT94y0Qnc42F3w6hH+iVfFpZaCRxUuiVmAfFuPxk+jY8WdYevmcAzxu2k0w1
tF0aSeZZmbYWZ6gDomBdUvwSo885dmZWSjVziZWzREKkhyZwaf4DSC3SmikDHP/iNwCyxHqHDLdQ
wZWX1htfaL5c0hR2CV1ETnfduw1/fZAPFA/xIYi4tN9WgUZnbb+Bk9v7/G9m6rDrvUvQX30OOjij
S3elpG6PMONfB974Vx1yhGTVcRLd1M9SqgbiO4ypPiE6QEUyOk3mbMAGtCPS9mvJ/uZ65p2o12iB
yb5P0+bLL3G8GtCkwMdwR1wAzDrJRdbL+xPkDxO2MbcReueIFEY8bqHcFj9ghmHYSwdtYiwIRgZZ
WXkFd45ayXyVuMBEj/XjKFIU6xIIYfrdYN1pSbfOkWsDZ5nIEGHqQBZ/+MuX5tVkcqk/j/M/jYjv
VD6kcy2T/yUe2Icy8POl3uJoAuxkBzN5fzXXC8AaxEKKqR0N63ulj/TJYSIFRqm2kpT8EidQr5iA
VPJAvlSmRTkBh0eWlWc8TCXKkteltFDgvQNEsW2WOZvseMEeVln+majpM/lqr9KA5YkKxR9g75/9
8G7ubAMc3FO+V+zA9NG1/c/IVhHf1kZUF/raT4WbDo8f/0PiDLxUMCw9EKySgFmMgbBStWUA+L5F
u1LMW9ofI7HrilBKHB+iFy5hmvlESGOvk27ZkCVdGeWU/eX1QbZIY8KBo44c02U3xiBTQFF/XMED
106LbvTFrVIcVJaSQRtDM01ksarUnPivXFw54M0h33o2bUeHIVJut2foPRHEh3M5DkTwh2aOrK3L
atb281lqp1oar+n+2AOdjDF8EZQyyn6NLHoZBa0RVPP4vxkptaDdlH1ShgNMylmK3sXMibj0dw31
R0UDgZj8Z98QfuDmSlOAov1xFP1paoVMNS5l5K84KaQ96HKEjQujwazq2C9EK5Lw2b/QhKGeA8sx
lM0eH2zERRzoa0wqfSyoiB9nze10f1Sm0YGo2Ydb4NxqEd36oogI0Bj01rnRZl+VSGK05Rvalz3r
YBj++LM01YAWhtxivjJvguqOkb3cIk02vsh0Tim4TVaqHYFi1EJKoC+1gqkvoj34UjFGuRV60J1A
E8i4KWV5dTXxVDqVe+Yqd5h9NA24EBF/7I/eYt1TVB/TpwBQZq+lvVDcKmpOleNDhpWM4DtpMxkC
wowXxYaJzW4gQ2RXzZ0t/Y9zM0lI+y6lzE2ZFmjIMxdGLN760xiVoLodgogjQmTzEn8OMOCywa/1
96tud1JDR22f9McDf1ES8DDcxWma9NAtd9CFLsC0e08qL5pROe0FsDbkQIqDB4W5Pm0hY2ETOoZf
uUsY4V9bScgPHMq8WWBS3pMKAX38qNUylekGRqEsLtNl6kWkxeC9ogMx0KnTWm2QFe5+bhSbbcdQ
R11/sFmSY3xbGjRcnZr/BhZQt43yZu73TQdBLfe5STmoCGODH8wKNp9mlbxiPnX69DY3l53+BiJs
AWGCKyBM3VcQI+PRLmqwhxnVzKGuOIQ1AwJDxzfmkqfr7MWpKysSf5TWow+oVuY2J4uAkM9x1hkL
xKqp/4t+yJDTDAGCvTu6R5iE5VlHphgHSuy4nlmDvyggm8+8/XYoJVIr1vHmDFsKZpZ83QED6z7V
JASlzYCHXVxCQft41shqD6JzVVu++7jKZT37z8dHSAjAdKRxBzwN3a5hdY/5fNPzjVnKdSVFxvrr
6jMo8G6cattlxVnN/BNW2N/AHeqo+jhA+0R64yDR7lx3y/QQqNWY7bFhnrdYY1d40udODuQBWA1l
o7d8okRgc6sAfSJTG8RuUpfHepDcsUEArPDWgHHuoJe69ZUzSE319hcu0MqkPXTkKX07tP+pgsLk
r1RWG4Yi6Xe3riuWvJUz7Q+hGi6GaGpBT1puA+y0hiZQRNM2JH+7vbdRAUGBjUfRSxnC6mbFe5cG
/Xkm4eFSRObgQ47FHtGt2F0gI+nKqfGLpGtrDEXvHpqlEJ5I0kfVbOQRULjrYrsrYOEiriBkMv4u
EHVAKUoOadD7sUMc+bsbNUUU+DpVLzahMNpeXJVEyuZQ4f5IFQGXl+T+cgtEZxPo7YL76Bd/GnPN
Dln/q/PJ+DlIVTlGDquVki3yF1I1DOOg7L6LwPQWLOOIJpKbROq8vxNObTDbAWQTmHRmjL7T8qOr
aOPHPOWd8gep3BZy2gqZrwu+cmGSXm1/JMqciOirlITSkmUZr3OPNedKT6GnBtHPDjGBIfhqUOlE
2PS9qIDFyXgfVMP7FJA5cF7mC9PLDsOnZWenXbykV2HNaplokAdk7uT9ukqxy8Do4J1rfT7HOlRO
20nuDgRm9rmw3Yt3hlELZrt3VlWRLP8tMjby39QLbh6GbOfxOK0Zc5ZMLeu260LvhV7VBy/aMqeq
jSkMbsOg4lCooAvhCRh2eGGBeijIIVxbA4K6Nqq+Ba113oPgXsi9gRhRWv7ED7V12RZq2h9uLOwY
4FO+bUQUoZ7OkZ9cfe3pYtW4pFW7Y0SidW2ZmIfsbgmh7qracRl4MjrLZoWskVwJfy5Y3zmTZdo9
I7OWAPNPJuJ4oL1Afj7SR45KyYKavl0Ef8SskOcA+BgoHxtTUgCfgK7/8cckjzFIrJ935UXyM07x
FBba6lDfCO7YK6F+zVtD//e9ehNldC8zHjNGDh11fO8W+WO7zx62m7MEkkGJQl6D5LfwcDGRjb0H
Jq6AXIg4tDrj8Upl9KH0QArcmJM672/n2rXDzm24QJiAWPr2VjsTBiR4qM/J4276m8iVJr59GwJJ
3+1/FHCpJhWzmARBy8M78MwF/gv4pAKJPzB/NLxAXTIketoFezPgom++mRbg2rbiBJBMOggsfIO6
Zy7crnTzToLVSEkgwCTgJ2IQnDcf8DA30OlegSfIe3z+uZjSKMqgJPeosMNOq94/kfN2Fss1BNBb
jCJfMNoRi9358vPERdMvCIENp5lYe4XOgZC/d6Q2H2vJJNgeihJIIbS/4kCFkxOwhRwekTqeLG03
gKZBtEA9pNc14ugeTs6fGZmDB5BFNoeHRNO4cWQYLKVtm4B4g66NLYsekQPV0byzswOeRf8zOpoB
VLyYqHanZ94V2ySy7nwbNDw7Z6PWMD/TqZgnx+SpH5CFI0WVSbnmQgqJniXUbcm3M/YLNxGotfuP
ANFe1dftnSaUr9SdU2uFA9GhR76vC7eGs8Uw+AA5XHVOE9bI1hjhi/nR/iQcXuOEMKL/R5ueLx4+
jaKtUvYDs5e0drk0erGNK/Jt2x7xGV+vYGDjJhH79kziMHnWIdmsy1Xjwy13tu01TF11m9OUy3KX
yCOODUakDzmpRVFex6I39Ba2yKmMmEt6kc5Hsqy6kdLm+3Dh/DPu9+qPIYE7TIjigS6O93lUrmcP
XN5QWQFZFhdu3zJntdkWvcyC0crOJmZXfgF6fQ2m1h+gEXlNcxCivVVmU0PKMm9n1qgCeRUJWHb6
93L8DKHu3fnSDeHWafHrR96mRuRm9Na6dcfMYReTznAmWNvDxtxI0fowX9YYFC7wwLLuKq39UEW9
H0AJ5PDUn09cM1chOIpoLjSiy16EMSyODNB4QkD6SWpjURXOGZli6H/e9McQz8mWwmsz6lt6Lgq5
QU5/9fidxAoLog3UM6gczzB3Gro7pbfQfJljJEMwXicTV+vxBymfu20VNMt7Ve4Hm9th9OxpiJuH
KADC78ZvG1j5tIY36TwJHWUevxqmeoedT+0N5qurlzfR670N3JmTjWuv86x0jhyyN0UfzbUgveWX
kB15EWtlL/HnoQh3T7cLWrFjVARwLS8ttwfjLsQzX05Hh4fX9TZYB5jZ4EULk78BQpeYDadXR/gt
tk8Fwmma074a/05HdIM3Ag9Abwn3s4eY2yBC7JD2kkLtn/50hXLC3dVxEqJQXUsEfng2/fvB7YPu
J82FC/YpXhaSwgKWVn+65FgsU3H+owjjwcETM4YdvIhsPiHq0iJ3hp5BafOCrYnVoWlGB9OWHwQP
/Ng3w3L74jwNmXzsfH1Nkh6oBeWb6He89rL/WKw7y0yMiRLeUQhmCL5C3U0mkvsMIf8JrjNekjIT
EKSBqDQZ0Y36mGYBS+dwYKC0YlH+fKUmpULsEm4hNYsg0IHsHolM7q6a6gvqtyCKEoo4I0BMIeMc
FQYC2DMj3dQ7GWWKWg9fSluVP2x4LOlnO5mGrqOD/XvgTSu2QMkM3GMM/KOXkoT0r87mEWqoeLiu
3SZ7RJYylyYakKn62zjv4gfwEPmAk76LcKeP+9i7Fuvc4cVUYO90gupvnklraEUSeaeF1ABeouOS
mKnYa4btRTidLofcTE0dp+uEgq9vawCtpgmq3OdDDtuLX67Vpuyh41F9Q8EU6G7ImdMIVH04qRqL
uwxzok0tkKoLX2+PLviHMmYp/5NZL8BLdHLQDpnOo/C9kabu3PbwFrT/KsPPrAq1+rdH1rEO1tnI
qu/wQJ2A5/3CBbRxWCRZchMhOHJa33BblWa3u71QHfYu955BM7BRMOkKgTK/FlKydwyiPPZxF8t6
i953mzesix+zs9IjvAKglxd/ZE+SYM41VMD9USiau/G6fnkGAW5C+jR+YnsmdUbZa6yfoadHGMa7
CXExYr/JBfjW8MaORSmzNas45ju9H6yGj7/a3xwuuQW84ujS2lkqlx3mWVilFTb2tg1VSeIP9w3b
CqyoZJxwZWxYYDozo9P2aOVdgkWhBuRFJ0G/Cw685yf/+j1Y5rGulHBMQVEZxovw0VIhSBITlO+7
ZFmR7vBEkKzx9kAmFSZsvFJymiQB0qZIdpM9NT1KxM4ZOHLAoajvV3WuCIdRofgJombWFXxhtm1E
vM0T+0IVxiEzMCwqaM/dleImUgl8opYka49jcQjHuJYQVWvZ6RQYq/BEmicvw7+/5rZtck+usZlM
X3cgG+6Zp4vvOs0n4TBE8I+0haHOV55sKqUD3Emwj/H3vP72a0haIY/wQQkC0mwRQoQtJiK7J8jt
za+iHHrpbTf2NUUgWxUy8e8Ue1DrvXSWrH2LKuL0YzwbJc3wasiR9tq3a1zZ4oOMMNgJkvp7C5ca
j1LQtdG1CL2gZlaaYTYzgbB0iI7r8Jvpvt3BSenGIBf2U+fr4clzLh1oL0vm32z7DiV5zZlUHxH3
MjWExopFM/qTWqHmOZJGsf+yJLyndPHf+Mzip3vgFaIkpI+50+tX7AOvvqvNLTX/KYjj7EwhJJET
dQAJ7+mVCfZ/tMt2EX2svA8r7nQk0zWt7UOWWkCfRSsEubagqjGBeBQnEtgyQ3rqk+q4LwNC3LJc
coQFmew3aHy+0sNXzPs0TVtZcnuLYhxFSzLR0P2ha7MTOBxWrK05za3fLbILXPYD57aBGeLRBH18
uN5DHz+hAfwtA0LgTKQ1ar+7u76Tj2MviizIkicppjU0FHVtf+1XwQRhBhEcQKWaJ/Se+z6hka3m
ywjBPfXX8zox7Ba9g0B8ct8bvH2SvWTCsYflS3sE3U0DsCHmhu3uTLs5YULbfjoFwIfj7n5773JP
ti63V7WG6LwfNgKSUfQbnaLAFRfzZ5PNPfxmPvqf+1VSun4ciZz3UxzzMp/sRf3SXcu7L6v6nMTU
EGmoBw67Gz7BlVsrN1rjGTMNAWEFwqcXykbGbDJPbnuDIcotjvdBJJ6w/xUFlck09j1STXeEoHwW
CYaUixqZn+7GXeh+EhFkHWZ0zDeF50bRFt/FK4X7KB035XmPbsnMMKgXtd+fVyPozkUJ9zxZefSe
4vCaYgUb8907HvyEHCGvdmqX1F4tqG72GjyvmYN03zpji9F0BqYFiBD4xUhK4QkTrZBygYKPEsrV
33Ohay1kJkGnE4SGiaM8/RpO9GMwCThj/pI+hSZ4WTKOoyf/8AIDWK1cTJ1An96R2vRXGv+PJpWo
BUxnSnC18rUi22PKC205mS7wSt0Se8WnT+6WK27kEgOKNf7JgN5zSZJ/WXjxE9WpvGUVulorBYiL
55IxcuEAs9vI5zfDUafdEVMXnl+cnGiLdiy3djr1khyFZsi7LrugjsBqUHtmmvU7hx0sb6dkfvy0
27/kMWmJTwSoEMelwvozVdPSPNhnooWCBtpV/jzF3ATRyCTJ8FY0HqFj1GUf/PVzJbmxQwfC1cim
NQw7HtMk3oHbtWerPQKHaP4E78zGFCr6E1CT5qcHmVTyZTw3c9vgVN6w5hzZpYcu1HcKZt0LQoZ9
NL706j3T9cfYo9nDlJkKd6OVoI1tw+Zcd2TmjQwnoJkMaswwJmzEo2Wem35telVpbXk9ev++5EmU
1+u6uCcwmtRVwKhMUyCMsZdLNvDX+35L/XH8Ntq0CITHAVuYWhie+KJMFhtb4gTpbgzoWPXpzz+e
zjSG/zkhRjELsnqeMgSWTAjLyDMjvPGKp7vhGMd8JRhvXqPLdkzGt3FJKv2P7vgV0plYTrDdaai6
5QyZwMoe7iH8nJfZlMk/V2KRC/HA/1Ct+TmVgeY8XBay7R8QODQrsBwv7InvbrsdnJSYPt1VilPE
hdkxXMd9tOajGvgiW7qqKLgvrhzmvAzEWNlPXp1T6aHtw6309pstJnrCVEUcN0oHwbnqtFx+DnZ6
48oCTXwjZlB+uuqOZOTH5uPjwwjwJpF8IVMYbF1RdGjHN8IPFM4RjiMb+ujF1uuJnyfJTHKeUUaJ
B+S/b5eBXtkuidQIoMuk9yve9pUDLkmcBSUv9yjR1QqxvoBj6q5puNUuiE5EVv1FOGPCbEi1V9Xw
BodLvNewH35KwWMlHif5q3EncjgJhnx2O7Z8SYNDBLhCaxszd8raVgiGMomqzj+yqm/rBpI4PbDt
NF9cWnB6e22fx1ju4ZXbJe2tMvI/7smvLj6izEjUwk8twwogE4yqu2U/A1E6RF/xvIG8KovsSLwR
UNlVFWpy3QtTYL4xtFhaqyLX51u8KDXzBB6P4gl7WGa2rIWNGPwYevhyXH1E7h60GIQJnbdsI1I9
i//l+YHXsIlL0BHef1LPhbeYcWPgRmOdQ/NIYis89Om/t48O29ejAY0uSYJ5p4ODauguh9lQ9ijt
2gBrTq/MJXqDX1HEHSdm0kQQbkbhIKo/glmFOa3YCaqHrxBf9J1meZrTHw97oC+ZLUnfuvo/pP4w
kInVOP6idmVy+pH94NVDnlv4NI7DdhM7z7DbJR5bIGvwzTO0YpZ9oYiTPH9gZT/x6qjWz9RPJxbF
UBNflri7cMKt6HVIy636oSJFye3R65Jdt0Gf7uDEu4FU5u1RU5OGx3DEfExtKnnrLPtv7jO2ZHka
u165ovSkxFEG7Lmtqnhi8ek4I4dwvdWCY1Zo4GgZD6D2Wr5I+HeIekPbaMAzI1g5B2BuI24LK/sQ
M2+VwjM/tDlBnIPVeJX1mEclYwaC5s3ybjr5XCSIIErZu1qx5Er+hv8yXznVUIt498PxD2v+ZpuJ
0liWKzE9CX1DKoDjo2UsXQjXt9myi9Oth1fN/ESbCZ11DoBxouKWJcu1jCMbY1ry/itevRfymEa2
z5VauOBjbAvn3zMoiUkfA4rb2RAXRXD9OLcXKQ66UCzX3M5v6KeED7EYtScdFQSyUpQGnzx7znzx
IFcTv7yjOJlbNdtKn6dIMzLRzZfYT8k2jwgRLThEiOrzr8Sn8l12rtkvXCLbVOsKhwUHELVxqOwS
OTksuVbAyebZ+BVWmVxR5/nzjD0LqBuYLA4LODcwzsC1oQxlC2RIsDmFWIiAfKDp6peLxyEvDImV
qUSYhhIYFSkA+zI9vxzrAaZz77Z2FcozT4I326eR7gHeRueACBfkmzX+xbcqswp0lsIHoHfkIzbb
YjmSAdb2Q6TYdCGaYc5eh8VUBw4Jz3VW4NOQT89u8juAXhvMidrM9GN3ITrg0C7TSSRyLdsFZBCF
DYbhW6X5eV9DA3ctbcscaIMLtQZDm8LeRxfwhOmOWhci7F6bH2q4RZ4LXfn6tk80uUUxOFb+e+Ud
0xRMMQssG+878Nicsnp26Zpsu20/xbale+FErtPo9uTZhaHIQ6l/rj2kzer57L1/vIwFGAShEJT8
YeochHkh99cttlK7lWwyammvTCJ93cDeZILxKTxeSYKO7cN1ym9ept7yXBn+5pFGhQ9hJ3tGsbKj
Nie8/cDRf6JhLuj2VxFRSdrfl2SGaCq3F6LzJDjQOK2sFR0M8Op4yDDzY4ikmQAzLz9OI6UpgBbQ
YznD1GmypSCTDMqEGUzppmbqfZ6c2sKRKeBQzPDzPeBuG7b+EyuzSr8fXfg8/Lvon1b/h7O9jRz/
KwbBjz9MFRJ95Oc8NHUSqeTNEwlAE4zRQDdNk8co4C+vPLsC8LvFbZjbYjIPQprNzd9yfFJa7c6N
hn3PYGDw7DNjsJOJv/hN5FOI8cD/iiaJkAOgjVU+Eb7BJuh47rOL6gp527PEnad7sast/xzgHvyl
/AEIpVtFb9dwMh9zti/YCeJMcdtUdG/gZ4G1pssyjooN9OEiT4gd2DcwsN+qKeoghJO1hWYcYxbU
J9Ak6V7JDV9GTX+L4qVfMC3Jn86/a5KrBv3yiRfS6PWSw9eEvR784D/lKTbrtuu6iGjLYCmTJmAI
gjw85T9y22oi0bTXvd0RE3xOgkEdW7njSRiy5EnLXYZXgAxDXVjj9wgi3IC8ogX9THeqn/j9nSXh
2E/Xe0FAP1TzMowmtKhYWaPGfTirpWmgLEgZPV64pHccLTxqw9Spl5dCOKjVYRwGXRawVKV5xqWc
uuGH1116+Y2SDORwlxDE6IHPA/cOg1IucAM4dDPVg/gBD5D1fGdF8G0OYvS+wFnugh1CoCj3iIUp
39yZRxys05TnQxXETS3J5B6RZRP7bSQDBho2k0910wXEtBzdKDb/leHSGlK4BHAijSpPCm7yVm0H
J6+hLjCmhxTjTAufv0aDskfA6kYpRKgMKIw1BIF3nMMYqExqtYX/RXxXrXwp7glZrE1fLYY6LPAX
/8IGmQNxT3zP3PYIfWVe/ZAOf94UfD8aO3M+QwIfg4mzkC/wSDxP9qFNTZz16jlLc5eHn5+2NU3N
ZCowrEDDD1/4XgIOW8gc5ZQhOIGR1cgMVnwTA9ch6gGJB5c2bWZUjvLvp6xQHg6CsC7UuajFBV55
Rz03dbPwsYeDDzRPThzYbJRb1jT0KyULz/eFLFivHk4yh1D/Q2MMlWrClxyfxajxRx39yaekACmH
KYAcbblMeZr7TVAXdvJ99r+RBDfH3TWl0FWFVK2O4k00F0iyL1xRvEuu+anhNJn1+TGqqSL67V7E
sKDBttgRLd6BSn34RlxW4gxL5NIwrZyR0GHpNJi6Zaqn3+j2MKORXwSnU+eeQY++X12xFgUfzWdE
CCrfQORs5lO9m1LawoQLcDzkgeA3zn4WWNBotAw1C7HH5DQMyl2+wi164ilyo4AkKjABhNZKEsgI
KkB2JvdJRMC274F2RNEeyBt/lN4bKGXFz22zUWzX25QCb2YudZ5qdgNuBHFETBzp0SbxmZQpVXey
i47dCzJpSIOeygzZ40fUts9aQIkCrI/LE+bOzk9gjdKI1HJc+v+VWlXF6/G32TgMwTRByHxi2bLI
bOtwLcezuillnAMBNGgLYGk7Ucevprebvlzqg6974eKXdVyio2/gwKbtBdzG7614tAMX47rlS7RS
udkpj9yXZV/020PUFKxirbAmhwF8Iee2NxY2mBKx5fqpwgnUvDwrnYEnvy6wpWUlFzh3OeA6F2X/
T11C60Vixe80n0offbTqpsMTHJzYykTPocdgtvuZT7e1OH3thRt7Gp5R6c43+r7oHC92wdPj+eLL
sNgBDUTaIIuyGRnLFzN0XhAdoP+a00PPdhBFlEcM3tYt/16pnlnyv9hqE/HXqwwfotILrFfpN/yb
Ha+yxlAX8e0LJCxU13I0xsBRf3z+69ymaHhRmGuomTH1DDACG26Z3RbPeDwbRpwnNs2P5FU8Zcjc
eeW7dkWH3aVml7v3oeOemx929ee4v2D7wBim6NSLhiSyuGNYp7yE28VUlsyK1r0zD+TuNeQZNER8
jLPiQAY8Hdazy8FjUsGXib3Xmzg8YbHKD9cFKiBR4tRZq8FHY2d82QDGuFWd1q8l1FYqMce8xvdB
PAX/iAkwHI2LSiB0dq0lJcM17tRQvWnh8u5cXw9NsTVkmTcNOusbHqdDbFlXM6DHrKaxXncd+DMd
ZD83zu4CAMOI+5DwJmqeqTwIoE1hSTPf0eZ1YicWKGLpbXmjjwgKzlGR5nDLEZRLDAdFel4q6dN7
tWdF3aUVQxj7yIc3tdFPMKW63MEFn4SnZw6QEaJOqc/jw48iwYiUVAHOIv19yPNheGK6ltC4aHkU
7i50nnx+rVB7yL0njYhwVXsO3ClfRS0kW3dEM0dI3umahXIYsjzBgAFS2q20bo9vLITtR7Qj5HFB
Y5DCuRYVpUZhFT4XB7bA9cmla/NrlY/CgqGJiKG9K5ZG/ytG2UEJ4nvMj3O+RBiAvl37bwd7dc9y
kX01R7wFeZZ8biidu5uLfKbbEKEaqrLaEKrqUa+7Gjkw62zT/BTC3c5hnmHBdfMNCTWbqIfLiURl
XAMLpnd5dbRLhA2LaJt6GnwSCXvs/YJQD89WqPOPa3JLZU2/h7UFubbHn+bBEv+rokhTKCquf8Vz
cJA0ttUiC7TS7y38HwkSl0k1LcwqkIfnbi6XeyT0UxxiBMSquqAawGsto9oLEt8JudBvrDxcgn/5
1Uk9WlSSlNo0cv3bZNcHg6DX5OfYUl0ruEU++URX3Zonv22jOx97ISSf/xn+ZSxCjqdSaBuHciQu
dG9ev/0/7UEWyOcBgm9UHT6htRfy0S8SFTCHCyfcy3r04iNmDno8NkOtAFeFyU90AloBExhunu5I
jxW3UJKzfNNWogIgE3QdZojkeIZpvTDuGprVBpnRzKwrNY2WBCnwM9GaUFH25++vgQA6g+1NbfIN
mUKqRHkf5Q0JTz5TYCD9tqOYVmYBUazxJqNuulkhxI0pak+n/L1RKkL/PGdH1WoTaJeurNmdGrDQ
hHTH7EMYcQLu6jMU4222O4shN7bUe1NMHULblHanop3tunYJHkIrxMiQ7xNG8f6vgYWKnqLNGVRD
t7KLwctaME7C94zRP0cIsbaOQU6/D4CiCITERiPDZUAyEuGLlGEdE15CF38dUKuO6kOquFyDPBxn
GdqtDT5wfRIAClH4UGFoLmjdVeFLiQEqLyYiMoJZT/6Ymfhsw/RASTqTUvmA9t8mAiP4uSzS3ufi
INvXgkbx4YTUcTzs4wdbe6R4zaTuVi8XnGVRW0VjVMp1jlhiKLf+lVxl7wX6Idj90yuM1hb+0NhR
15WA3GuefLb8vYHd/BCb/Acgr69DhXqxxo7wGWXX6RByfsUk7nNykKxVfLXD3XJWPEjWhLGeBGcj
wXZAfso1VkWWLukuAs3WJbKQrae9zfNWK/ixxpjPOU4KVKbSeht3nBtK6KxuU8u7SlFtPZJl3WOF
Kpjxb/KlOGK7cGXuZFqy0VRvLfpYsZ4Tyr5MjqG75hArm37e0Zp/n9l1LMWtfO6GU+S48YL3QvGP
ZwdsWWWTe8SdaZPbidxAi/0wUbhOYgYAS7/t/LR8blDS8WiLvfXXirRu04EDYTjLJLZKpsN/jret
Ua36wdiK0tF4xtVzU0IdUFlxAtITwdFSCRDI0VqLcX2+fNK0k9l+YHjPsKVTZ9QH/KLZE68qquaK
zskLbGhLzVjZNmk7GpeDzTWoTGN6Y31zAghjw1nKyIex2S3ocYbkyHZmpSwmLYl6CdipNVt2p9NV
9NS4tdpEjYWrN+TJOjYGV9SUCL+CxNglkdnefz36fZg3IHvBA/aBH/UX2rC8AKwMHjrEEcPNErrk
jUkPJQUgcCod+6H+MpNVye8kFw5HNLjK4J3ZkN8FuAXtj3/uuj3w0LundGjXjpDVsm9DJltlg+fr
0grqhTqDh71MLxJWDPkTZVc5kqOrJiuKJwJuGXr9irWiNyz6s1BpI1eL8jiydWAniTZVTTzYZl0G
EffpJWgnkgGZuRJZrOJbpJ6L7QaPWjPBKiMSN8TCevZu+pF/zKpIdpIu0DJxAXK+xFJYFdIXaZr0
faj1ARP5uiwDzlTeG5yb9DNSYND3IVUOWZm6ctn+KnYXn2rLIs2vNuNNFk574MmYAmTeW7t90+M3
wV0OOXQSGNyv8zWbIz3TiLn5iAPUwv9moOGORnzP+3UJBD4HH+IQzCeKF4Hcso9uD5tvcLmEQyGt
rMhO8ssR1WMfN+8AAjZ0pQtUgO0ZhZMufPloiW2+nrEvICGBPgu2czGV6j1JgA7z9fyOOJUyAklk
NJbzt1bpxcp4L5jKo+jOcT5Lw+aG+Jaj8dyIVAc4AJiQVxnPz9Q+s/i22ITQVFzvpH8Kp+di667E
lmLYWSu7HFjrI8mOzT1MI/XwCp7l4dtUKb+3I2iuJE5YXOeO4aMGHUEraFC/UPy6cWmrnNz2qHNV
wLxik6Lx/ybry+x6O6sptwiTq59AeTvDC4dI0XC7sYHMQC5b94aJLwLeyh65BjIiNpT6WYNwJpdh
XGxL4mhCwI0TvA6ViTHOz8Ho6qTEHutIlLaH13nvweoAoEZ8u1QPBY8dpY7ZVqNBVQKIUqQi062+
sL6VdkFjBrDvNxLRzdfxHBOAD1PPmUgWjJ3iXW2kKgID3VCUdlcTdTUq1+7A42JjOVQPXSVXeemT
obcpHNaP8rsrbzba8RHa3sbZHRLh/wI+Mo1wBKrcFB1Es4EpHxQPTwtiVsjdychr30DoCtXoP586
pFr9VmFsNGHBCt2FligiW93ayNBrQJ/1df7j77Gcjh7c4Bk2hQOuSij0eKBiPftXGWEYgqByb6cP
prrPIeUwhvWVD5rVSy/QgIbiY4NjankrAT66ktIkFyIiiqz3t/3ndMbAwrA2MIcWZhNwSHwNmgO2
d4IEGhjn13Dku02P4pb9aPYaMRZnGQG6Z9w6fLVz/RuCfQmrYbKbUbA5Mm0OQDMYuXrppJV0+rs0
3fcAENidpaDU4Z5D9vjXCL/EF1089aS0qAc+GX/6Pv/Fhyfiwgi5AZlM9asKIa8riY0/t3IrkiGC
P6xVwhqRfB1++Ap4sdIl0DZdDkMqggDhayPY11XKsgNO643unHBnoQSxuZv+mySqdyBbFfOXyW28
OAFbq66MlwqWR3MORaTAfWHCblttQnLbPLLQ6WPdn9aejwe/idnU0dTLT75bSoFpa2IL6K1C27+M
vLQ1ud1EK6A9SMSwz4xv4dtz4iAJ2viRskTWPU/m3YkgjYeBJCmOIBe0+C6VIvpSy1eOjNbTWtgH
84uf2tBVdQPLNTz8HtnfQcRStVZK3Wcw6GaTEzJ/9ge1kL6D5gmJZayUF0UTOXewrhDoemfD5OfH
reZMnfUhTB0KV+rdWVonIy8YszmPaRAWTI/r0F69/gmeXWqL/cpJRsyR4WmyMw1fW1oVtPTnfXbm
R22m7lSYu/WubadK0dIqZlR9pt90Dy7B6qOvb+sXFzkUGAIxMXuaiRP3RiaHhtKeulaQA6cTNIvO
qD/1TtB6MEOvl2Vwp53XC59L9EW/9rzoQsG7VHGvKBgxr0GW0GwL3m4CwDhJ9dJELbefgj0cEk9o
HUmHqHtyob+KEEcuGnFaYlGol4hHVjIdCZqESW0BeSoQbN65Rq9FYh0tlz4H0LhLaI8PCx15eDHD
fSdcb9Xhocaw1B6ZHZcHFxtKo/ecu6vs4kV2RdLIiJZndyR/kUVnzgOHGkpQcXpI7SdAVk6jJoW1
jlfc8rw6wVi2HUVHO608jd3tmiCEGw3CmIBzejmmGGWlQBloJQwBWUcle9uf0l+K7xxazC/15S6r
vlHxMjCq3VygDAKsS16XBPLrphT/xoSDPLt29wLN9XMxqkrS0QAD0c0vslVQU0+T/CuF9vAx6r0P
0UFLiD4nHW9CHGiWMiOsIg0T/3DfIM57ZfC4m95+yKmieGWHANpkYcRLgbdTDjV5+e003qbONy5k
iM4xLW/bnImScbA0lWtj7q1QvfGXilmcQHb08r6zQjt7PO+vMP5/9N6z5P9lD0QZ0/Qw3VpgcIzo
Gzg7+Jtnd5FsECjRImQoxGfYfgrHgWoOxsYgOxKZeEjFmdmu27mO82WyeFRuHHkv1QO7KCH5cYZW
mpBJg7JrDzz82J5eRT/SdZl7D4XAofqqcfCQ3iLr3Bw/uhJuXfxoAiM+dePnU+ECEM23YiVuVbZA
slDPjJDdkSjc0+hmdFup9kFzRd861+rQxFqhHb5XAYiTbFLIhDUkFLOAWQIydgVweqi3aBfWdefb
T+FNFcFbYRT8qGNqfhr7/RLUDAd5MUjPHFmF+lgWjz90G+Xlg0FUNL2GqasoVeRiWvC9aOBGvAdi
cCKKw5QToPATUGJ89x9Jdyzs+h2SoAYrBsZrQtySmqATybZUl7byzcadqmyvyfGqjFE+3zjzQYot
aqE8GWkRvbV9/D9rq5UIunmhxZt0iRuepD4JlEd6jXno/tyZqUwl+Jnoi5IfMpPTMkZOe/Yh7jZc
8Wqd2Q+6HjijpQ+8kYqrUpGF8VgEVM5skBzJ1uImOKXwlfIm9Xz4J7S1KmCe1+6f3ma7AUB4qMsu
Ul75SCq7y8Cx0Wdq8/MTFFty6mmcjS+wVkslfHUDoUgpgUlmc8FOpjli+JlKVwXX9P4vOGKWPOkY
eMs+NmT4MkNSK6q8vw62WGsRMdNJ7Viptj862/glgqQy60gE20DG6wC0eczfLQQJHPCwkodeVDva
YHDkFLkOdmcRDLtVP3OEepfU+Mr0Cs+xgjnVjBMAVAyTXH1s6yRG0opZDrRCIeEyNrGpHOwzXBqJ
QCLpJ9AcD7LE9xTd7/pOhUVfvg8VHzr4ETCrSavBG6A89bK5XWysQIU27qemGoF06imNp2LTU+Ew
l5IPuklWj7SBryusFQqgNIK94adgkZUU2qwtKaYZBCqHnIf+KVEPYK/yVeR/AM9HvJFe8/4xx5qf
bYVtVYTB+JG0oCwUfn7vbF4afhxQ+5261C71w4RhSfHiikhAw7eY4hXxEuXU+Ka98kx71r47dkwN
qC+HAqKBRzfz4GULmMLdGnKIEwdVoNUMzC7A58FCkD3SGtphB1K0nlRU+O6Ra1eCBnYT0plGtUJi
+6AnPG2RLsHAjTVjN45QQIEfPccPuxr4wG5lfjxCLsdHYQBxzotdueoIfORsaVvV7VS4hBvrlOY1
E46+oCdVxTgDFtFOqeLx1MghP7/zoRs/7DqgVYVML2VDfXlI99QcpIPu6jK5sBLUR2DkvrgmPiL9
ezRDQ/HMtXz8CXTkjhavVESnijmRwVLBrVvOktGZTOaL0CgQUb0OoCoC6ZhdlA7IqnU8LaiRYcF0
QGBzb1CVfSD7fRyhin+fazwRx5yGjWCqrmCsOflDTHNT3CXpYHCJCl3PMELmG3GBI5mrbt62L0Vs
ccV3lfsCnA9Sl5JTPG+Ab+TuhYjDgyHvFKbLGOITK91nxdjdrqhFV925aluMye814XvgEvtfVZ0i
de7IP5DI4AEbTxJ/Emh86kJ7vD/TDTevTPSfg+BmYMBhK1f1bkyz7u910FdFrOGxhNkENi+l/M8Y
e90jNAaUjLFn37L007gXMLzX0ocp6BdW1SwddMjrL1x9ystNnQtcTCfjNd9u3yElsNNeOYtYuqRe
TkzS2MDJceqR1DQ8IOFcTzs/VLLPiG727Z3r1H5l7FmOtQxEaOh6yT4wqz6ED2WQLTnGr957folm
QIGmLDWh7f6HN2CT1cGozVDzWVsGhKbkr/9NCLsdzFNevcnfdpdhOyNNpt/FvpG4aGLvfpBBkhqS
iozcvYZmmcGr3s2pzjOwx2Ozpd6ZNai9vdzk+08qDw3LkLUzGLt+9OoRNNCWwTM1WbZsfgJOHoBt
va/b2qKGKbbhUmWuf0mM0Mp+YEHpcPQyC/widUKrdLXZg1+LpQc3w3r2RMVJ7vD2mMGKKtTUHBCp
dlXlbSqWyE3uIthQfI1lue6UIbuuFW0ckHHP1AJRPDB+HfPCJLOA0aqb+63M7KK5m13YOebKxo8I
5knT3fKGf2MGUKZDG4O7jHi88twnxH2+a8Sz9mkckw64dyErHYFRAwKAIjotccI8ipDbWOLp+6Z2
iKtEUISqXgdrejox8ZZ7GF/1pWbl7WbkjbFfwLkgxgG9UMrGGPUyI51cnvdQmsIbPe+XFROfBk5y
Nz+kSp+MwiTQt71Ieb31AJhzbcN44BODCMBhqUEmgOLG9Y9FMFikANopOfRj/rnT7rn400+l9437
AXn6DuKR568xrt3wsq95W8dqhtlP+CczJIXeGb3VsZrxJSmx5t5W4FckDqPvR19tC+kqrgX31nst
oVYebWf4M5p9dNkMR080xltnwiR3a9o20vGquZ7iCAjfGpgOiiVm/OnlZ4X3dxRtMXCmbcDJMuip
Xb7yatAUkSzaw84X/sMu/F4vrj5mDiCpgyfz2YC9VKYezVBENCDJAV9IvJ+8OhrKBSt1jpl+hMI7
c9oITWJekxYJoJ2gXzVI2z42f8WQLytw4eXWa4nkjA36MQYJAQFRh4GSrAWn3heehRrP7fScBTzt
lKWYlaDqGMy3z5Q+oEi83t5Emc/ZIpGeyV/H75SNsNGnNkuGu3e+J+9B68W1qdl5BNtdWVBy2K3O
RFZ0TN0drj1qhMARW4aDwqugj7zmsFmrLuasycPs5L3YjwG27cdhl1+/58++IjQWQnM74yjg6VBt
LPkqxq7ptC4lUI2LFo052Ci+zQnUb8FaHr4O9ZEfPit6WIbTnylV/hCgkVcSFKXylPR/FWBU77cx
4mnj9NqSvcurkwlOhu5Xp8NiO8taoGzFmVRadqyHso6GR3ehBMnhfugXk0ZOGha4mY8ZOMMDmmfq
UuSMAe495BSsb2bn6vjk2o+/bg0JmoZKFtME9LOQCTbLzAnXPexqRTP+mcHAGZ+eh8YnDpJxYzJN
ScIN9L5Jl8rqxJmejc+eC7vFUhoCW5YL1y+HxoGz6Zaw7g+L1DYhDcUZhJNGnmytq5eN1VRe2e/E
5RPz6jTJo8ZyIlIsareQcK6akqtTh9nTfDxqOuLfSxWa2cXNC7shWsfXt79FubTGHZ9+uFZV+EY9
vhscETgtZ1FeBf/uY+zZ638lteRL52UHd2gNDARsbGoRrLAsfwYFeczS/9FQgNYhMWYo8525vFt1
9C0eilOrbPo8wSrCH0VXwbbu+HYIQspRYciYwcow0Jj5IDuF1kidR/2Rn3rZYQdQga1TxJae6nvX
JFIcpQXKYGOjRAYpsPdvzRReZf62H/8K0VuyKQ3VruiECs1pIt/NYZ0mjsoZYLxeahkQso8AbOXx
rP/iUQHXacpUGO0Y8oitcvQLPNeuf1NwAy5IFsUVKXyA3swOH40eUJJ9IO2XcpTtu4f/wdPO3C0o
zEhCsvOKZyGLps4/FJb3QLVkK6Ao7Xuq4n35YmJGxhe7wQ1jccI/os3++h51a41Rx5q3LVdJPX6C
PW4mKJ6T4EYhIDPQnc7ElZypZnHJMmJxHxq6iB0mZ8S7BDmG21k///7f/QbJ3B6lLnPEKl9FzkLK
EV91zxvzM3Lcv5SGEhzrD/Q6JYU3df5BO2mKPlVAoNuQOrddR9MIGpjboBrrimhmSDalpICTbzIL
5XDVgiCatpCPK5j9QdPtVOwAUGk7HPrRW7fByCLCRDdo0saoGwd8//lAS9A380fTBY6x8IoXCgR1
05Z6MotCv+dJ5B1e7hBajLH/cxPjwPI+2l0nBccgwOqTC9TECzlfC9cq4GAPS1Qf6Y5JumROC1Hg
A4BHaV/6NDVbbF+7D7npV2H3PKHGeQHtGzPCoKHF0Z8YSXpYTMPvO3X1Ow1DkTXSQIpl7cBTvbCw
jvhvTvbFL1+iWwjGaYoTHw5dps3Uf8qUc/6R+GeaOhJL4cfQJ2Lai6Y+M+tsTumK96LLlRpfxSNd
JXieXidXlWFNucmZ/6cJHxy/h/wDloz1A7rK4Oah+vwfJF0spraT6U6C5AV2uB1pyZqkspoZ6sGb
4gfJ8OTzANr2f7dzrVEUp85++aCyyYrqyvsvP7F2AKQN/EN34thCxDTuvFp7nd6qs3Hl9HXwF6HX
eNA5y4OVrxIldmUbr1jHz0Z5FYW401WiS5U5vNELzPCagL5MLVW3blxUKALa5PWuycwd1UQtdXhf
huQJ4Z8LMwrr5em6RoIMI+4KsqRgxCU5EzSjzJ8wga+rYmyztlwWLVAe71hqZxfqk4tK0kUEb7SM
H7gX+0N23H+OxLL4QVEGTk0b/MEtYfjKPwkgUKWBZSfjh9gXOQkEAAeY/IoW9rj3tfR3NpUQJ43l
Bdk8G1vO3dRAX3zjH/zJ+75N7Gr3QKykMZLDaGzGC2hdpJ72Mt32BgV5x72sC9TL9h3N13fm+Wjl
NgfQesA9yReKQOqRF/HK6s2jqeCsbXKubkHHtczbU1eEKCgdLxK49pjIgT9JtY8v1ujs7RiObM68
RHJPQgo2dxSEQ1lqt3KCmMqe1xON+2k0wSIgMflhYVNsCiL4mpzQC9/CnrfNPJMS/5f6c8x7WqLy
6sY39xPGRjkYMjDmJbfLSMnWXrcrTGm1gOaRq50zj7oHXex6lbHqoMU3p/SukQbr+qsZyky4JpfQ
FjyXc8YxK3grNU+pLoPCxz6bXEOEofCDESaQFFViFHbjgQGM75ok15x/BHc5SOhrzTY3gIlSyzzi
pJ5ZsbQnKy3/2dd0GTNQ9Li13p266nV1TzLtFeKv4sUY9VyciinEl27AltnJfcDrow3wweuvpQru
sqLAaJ1/p14V2PbDv9B7FTgyQHV5pUu/N/F8Zq2QLm+8mGesZSo0K4qrc/yvV5IVvQsqHCv+AlGx
URIjmEDQfzqD98z8q0+AI+3/zTbxAVYk7cEll4loFWlrWlGm59aGsEob0nU3ERZfIgW3CWenOHC+
n6x1Yb0eagFQCDYAjLLJAoETS4XcFpVQhfrxoT9ZrjoPr1Qa4h0u+JSZKfxl4GfxyzHZtX+DlHRH
n/wo0ZKbc/vHSswShCrJq514Od2RuB96A2rgWoHgK7MZXgy3GxwGqWUnK1rB3B7Lc2YQzjrjWAqQ
6ghT8iraxXh9xNC7yYibF/1RA2w1OrJLqaDWBsT5/k3fESv34YNa+UVx+Gsa6AnMRndhT75Emz5Q
nhrgQ4Zp71ezuR0aBALa6DHL1nHolI0bKL0reLcXWI5POpZ5TOVogqeaVLXB+X8vC79W03tDDwga
q8156kDvG6CWtd8GTl5JD/zi9oeqn+i2/9qKtwpJYXgki9cDxrQ3EQt6Ci63OnPWWbADPKRTbu9I
Ce8EoAXD+e4G+4ur6eIIiiMqBloEidBy7I3jRgywZi9ZCT3cvjSgemEm++1xYdVZD5cqS3w0hQtL
V+lQAmeb309JX2EJaydY53oulclCj/vvyiQ38LBCkROTzw/iVoKquPdxHiSJlKHkDnjXyxb4Ondu
d/oxBiTAz2sjuoql9GBvLNo7BpuPHg5hAI6SduvaAlSkZzGLyR2JdhSiNwPSy5cdSDQPNoT2L/Iz
mBt41hDlw9PiTeZbY3OXhkvAdi/b49Uk0fXxrL9rg69XweZjAP2K8NSgWAH338hMhIc2L0SzCTcF
KmbtyG4xhDfPh4nmEILfy/qGBDwbUZeZVW+Mb9t08jhN8kQ87LxsZBj6xbVzLJgOpODJnFsIzQti
+sBnXn3vPTKOwUJG4hm2KGBt5EwkmCMMeOtE/3q5/GbYBPqWRejOh65aPpZFB2iTkIZMbH7HvB/b
XQNTo33o/Qifl+vXNiOKwGOI5Sf0m4Wc97mVl0fHF6jTVxUG3s6UJzzkrb5A6hbOfr6ukkP0I2v/
uuAdAjyo01RLZfFlsnvFEBxtwU/LjOErz4es64ip1uNxCp7IM4bcQtFbEV+ixN/vNy2mrpS/TXAM
YPFLUPWiEQEHaIv8HPYb3y8oG8eDtpP1tRiY02QiTg2qRuitDqX4q7fd9131dgSqWeaZY5r/5Jnp
GfA3k1vEInyb0i+gR8r8noAKT87FR8rvahnQgd4OQcTJRx/njKx+4MRZ67Yol5y7k6/SFvCNEHUy
d5W8DJnP8J7EQVZJNkbPheKO7U9PxeXrr+o+3vCdcAEKYblpk7v4kByNcC2dfntaRrK2QyPMXTlF
G0uBwORZKYK8r3ylzSA6qU4GgXyyUL5dHYaaHvmjpWreu17mBj3M/2SUqmKZovvYnls3tVc2QeVV
CAH5NIr+DpUJ+OI8p6flNdWMy1B/Jz2H96YkLPcCu9EheDj6+vRA8zhMdm9D2qJuwXeq1KbLJtyi
MSGqYJpTIImwb1onXlf3VJT+u8jSMcJqmFWOuOyy6F0v9ecEFx3F6yNBaP29ZLjIglMuUZjQynDy
aQJ8MPuRCT9U7SmPD7+gWAkXRywoZ5ZkzoPuhpTbupDkMDZ5y6SAJ5FmZUcY/1y7L7EvZNddV6aa
xBNZxZa0G1mVT7uLQv4vVlDOE5HNZWMS74ViJkutm6/xmUyNgOGN5zQLpivwS+l5Uzo35ltZEVCF
BwqBbjyfsMBFTahDt4FRO9PR1H9a/px1kjo7zgHf1SJLlIxOY8qsnYfufeMsiJDyUtfLq76ArofL
KhRUWQv4jWqV2GRyVKBWgmFBnb4RlyXB3mFGNhrY3InMkNdFzkXnYyyfhs2zkxuY7gvKUYr/XkUA
O5qOsvLNSpN79koHrpCZrOgAB4jK2rdLgCnoitj1TXvxw6/hzCD0+PxNTsI4JDJBOADRBovL1oLr
PC7p3gIvhPc8UZOgrW9l0BXhp6l1bnCEbmb6YveVplgESVXrTeHm+2AkwHKfk3CfqDWW1OxgD96z
Tf5wvXrromqvYBQYcq4NQoBNC+VyasPFOfl7I6pWx3hwPm+voadk831q1tYl8O25SOuim4QDYXJl
ywMOVWox1/TX6DVFp2k4W1Ojxm/gdVKaa9HKIFeHebVyPTPZAm+P807/e0fEVXQh9+0enfoqk2lC
2xQzv2fBq17j799TXFKexa1FvhUap/OMRI5JFEJ3qJJtX2x1w/a2E7KTzCxZOsN2p/LflaiveEU+
QO0grCpMBzLx0AT8Fik2ZhfZqiZUsBIlHIzJ0u6psdeUBVQoJsVPYLQP5m5RW87x5dG4UdyvHETq
gBNohOpIGHHEUBV1Ek5gL6D8ySiWYMTEDv1RB72BUPmyUU81coNH7Ekcs2fd4Fl5Py4jOOfFyx6X
YO05Ubx3n2xFEU2ko6XCqDHJge7ILFhaJ5dHoVkAK2mbo8Khtp+0+nJnNaQr2VfznWN4YKXLEnmS
owxuVYy9O8yzMYgLL40sP8XdvGpzbkE1qE/Aekhv112ij6kGpF9AA9MHnOhnmLqloP6iS+Yfb73I
6/ShcfP5WoxFsBGmsp9DWFCPQV83HHEnVcZMJ7rtmLgLhVqR1fu8iiuewl5A2Hq00Hv/89jIkrJp
T6qcBLCfmJaKqdwb61Nlvr5+Um50rhxJtdV5/1Dp2eAY4QDOyry4NyDpH3pebyLuSNvAFt+bjnQq
kVMzRtbQxnU1ZW6MdH8psMSSz+eHuOxdZ9FwS3rYl8JRt6jKZ+RSyjNNm6ZK1OWJUyVoCuOvuI6s
rFnu9guasIutHr4JpLc6/M/CcSTL4cqlWzLxIFwTX/BB44OD8IO/PzZtSCHiKnY24l909Bnsz2/P
kbstv3aAA0qDCcewsVZLWHBmKFqehQ5TcxTl42KVVgG+8CJ0YRrbebOJPDjA2yzso4mCr8pLn4Au
1FoAQrwfJDbWoJG3QHMXcmMYYDQkhr9cJHyV2izHhVf+L0Q+AMSyfanKJVq2+XyclmpG6qm1uyU+
wIP+kFNoh1gPY37J5JbL+0eU17ZEd9fsoAiUTj9WvoDhE9MJF/AwDGDXKkoVRc2LEimQz2+pGFyl
rW5+LEvvN+lSCItafilgXw1By4if0//JvhaSUioIGqVM4NNcs8DdUdp6cZeug5KCXMPpR5DefnFc
N8pOqWKSMZNgtAM8rHzrqeHCNeOsjHEbzJ4ApkyMAShsgESPKlpNdtE+dNB9hlbvYF1v3vUwxLQ3
z3d+ZrK+jrd82slxVfx++4qIQT5RvxOV0EbpDqcyKZiZ8n9iCNOnr4/RjonYPHBlRb9KGhX1ZIqw
BZVwIBfa/7adrymXkeY7PKxA9qu6YOFoYABn3c7lqYoOjaKxsbikoCdohRJDh5McFHFc72RsuwLt
RUSeRpqpXkl9rBIQEOdabF7l/+xgQ3FEfI9ce7rcwJJvPtNSbhEKYISvk9BLqISe0439g2NefvR8
oqZ4NsTbAZJwRpwnsvbyfUyhDUPJ85yca4vkQphQL7OKrOFW94ocIX1dN6Rq5nuHS3ukJN3LJVg9
bcwsXuI2OzawiYyTcFiWiHSYFaBBtUy2MNbORS6wDSV0wJAhwbq9v1gNYpzsv25jW2tVrMlS4acF
mIyYZgark4kg2ugwyivrH1EKHZYanyiB6z54dUV83EJv76lLxl5RHqcnSOXSISpdDNvcFsdnjoHC
Yx9LGA+24pL8dQXoSp4mzfQ384EdWaLI4foBli/G/t+BZDmZ8B7ul5FBqVxIvth236hHy/jEDf5e
tMux4bDKv4SqKtC22fpimsIThD1b2CVPww8WQEYyCuG8NAPTFRbEYMRk3lYGyqpVdanYCRmL3Z4K
7eG9DwAcDBXCJQ720qH8i7Z0PkWaiRkDA63l2URMpWDon1Evb9ynOJviMJ25oB5/547mmt9ooxOL
3WEVgmGrTqS8nXMNHuqLeW/8k1vyY9mmIqUKQd4o59urdBVvM1WLSArc3WHcAsKj2zK1JF0o5c2x
88KdNKcxinbGyHJWEDca/whEGwBJcK3nCr29cm69bCFvNVyP4zWPneXwKcGUSh7lb7UgaQygcnbF
nIO7fa1SD8t5kE1C2Ntb66W58C0hVB3guUL6jb3/tsERidhho9aHtIRLCKDNlnBPHahkjSuZa6Vf
Htw91OyVGTGmN+lvSz6SV9Dtfxut2B/Ij53eH3Ow1zr/afO/KxjzRT54GOipo9xNeLy7xbzvxPQL
dx2a6TC11jV+bkAdHz60nvehPJBnXtmStyEHgvumz4nh3O2YAwVT0FOzuSQY+BWoKaql98DUZyV2
TyWy3aCH1fkwt641UoR2u7Mjs/QEOfZWuo7HqQ1pWIODqe5X/ewNv4xIdGEiv+IukZR36gb76VuJ
FEEv69HDfbgvwFkkmWCAlZkq4wovGpeeivfw6t6NMgEiNLm+tR4EpDNtJwYibwBCVP6//NrFYmsd
KLrFrH3VyibWraDWavDf+xsNTVyrOQyTbLXBtuJCfFAOIWkbQKkAW0EHMBrpENxjTi7FtHNJQN8o
+R/TkXiPvIj2jcvjXWGK3n5DdOOj32GPBIINbPkiLvEicDZg1RfJiOAWEaY1DcBquVanFb/WB4lg
Gf+DJkv6D0+3vPCWPYkf7H7iOVLXx2p6UrdSjB2M3O8wNrh2t0ibteAzHjE8k6Bod8zA2K+wHNB/
Fc/h5DLucJ+vMhaOacgDnhtrKDH7z4Expu1ztZunxp6NSHZdUqEOtqpweElmoHmI7Jv9ds22CsAW
D6tTL6JGcfvPv8h/7NTkiWdziypxpQSEdKw5sYy0ZCrlQUd8TT5zYaCQjDfw6TQ4xiNBdWBboZZ9
r5nrVDtFtxYcodC7fba9xQP5hlmE/eHLjluBUQbJ96ImZTeF3R/O8XeuPYVNzt5maCuw/jFf885d
t/NKx6k5W+fkIMCz/jTXwvUDE+ZZ1soYC103+siLr8hPSm30gO9OFsG9IwXjfTKlJ4qvHevghGNC
yGN3uyo/axAhw53JDjzNEI2eKWnJRoDVb2iUk6okW32cpv5i0RT3g14F2MyrXnJM/kqckXzyM3fW
iVRwU95MD3XSu6h7UZbADufC+ekzxk8IGqQGXGHJGDe77uGEuZny83X4pt/LQ2OW/+nqc7zcTvUe
+tZGvNeJL+dUqlMvOFXmxlBVmbKCDsa16zfciYYrQaMDigVurB1SeioFylXjkZ8P9a8ZsUfYETsB
Hdckv2z6q8ocJ3dWRO9WniJCGzpOksQcngnQkDGGC7WaCv3cD2oz7Z2Khcz64rDQ38cOF5S5jg5z
MWtshazblQuYiURYY9okSFOM5abzMxCtADxJniZBoz/7xo+ZgmIwYq2yJWmPxcuX1B4ztdteGr8D
KSWI35EAhyemsteT3CjiYKVPz8cnfHWAldDYuVgzA3/+CHAEEltKVc1JiLYMjE1eV8j8qj3HkRwJ
UbCD3FTmu2swGQm9nWknm/017mXsZbcabPT8bcOg/gPhnGgKA+A5Kk0QlfApchHnzeXkESMY0D6q
2SsQkd+8MJb1fLjNwlo86J+SjFzS1UZO+H6oWZSPX+l3XqtOZf82CI7qnK1A7jPVb4i1//O3NlvX
DLjCrBLo0jnRhzea1jOMpRL1ny0rLr/gye9TUrVO5IAKU2wADs9F+e1AS22Rs3ceaQNEljfsDuIc
+tbvndmJgl9eG9/1Luv4KNwv5A+Gz1j3KrjQu3Yqd42IrU8EdI3LGN3g2MO5tDYYLMOzMdB7ME6n
L75AN/X29ozXRer8iYG8w6nMRo0VU+xs/rg63v4QeK4XoO+SwQOoXrXHryd1KNQjDD5lXzOLtaqh
1kdC50ZM832Wm5hgLb0wz4MaXuxihN2HUeeW2BgqC8BmUqP3zUvwJXk9XTfWuENVgzCw7/PFcvu+
EUvgaE8p8TznKV7zDF2UX46a8ph/pF1B7qVt56gAvpppH5yRh4M3ajkFbBbn0hYO6g5Jj0wkZbr/
TgiDMNL0uE3qWt4XoimCtgZ7SfFGYiSFlaWpqfvALdpneVnvctA7dzr7oAtq8u4Uu0GZB4iCiuvk
cFv80t26CmgQe8ut/nJ2cvnAmX7DKoXD576w3W7mFkR0/UvdUDgbHGdARPR/tKHN4fdNio7vy1aB
yldNMP6dmgkrloq1BgzyjQXgRtD7NlOYaFU1sWhSIfVKZxd05CL7BiuVrFRta5fGLMOzyG3yzFjW
m5HwMkGToMbsQMeMo2MUmCnjBbLDAQyJ7/2sPcp/6Ul4iPTFu33UsMBcLkPqe635849RAbydgIa3
0UCnTT1ApglVqsALrqhsnH76KZ/oTyf2c/lw6HEnmBjIGTDBtZApWr4hzKnYBtOwH2NhKwgs7+2k
cMuzhaj3t1KhRmdNL//3f6ObcChPRfI70qowd4P2hwug4UZsPnLzZWyXzXSKGdGMjGNA5kAnoWT2
CM9v6gXMARq5Sod7m/rLwV2/tguV1EtWsqZH/QzYjYKFCRBcA9LP+a9KcOpBIT18B4gckUjPt5ms
DrIxvMzMPvnKHjvWQHCMlfi6EJwo/u2da9QadNpG+1Dq4LrQZPnjJ5qploNbcnDo9lZPo4kQlJ3f
CfkS8rbU01QM1fZAmiBm9foI5qkkQHd9UEXVxd8jq9Iqx1wwGkeOBkfIh2GfFi+hYpgjzjG/AaLQ
r3FdFCpPL9aXSkOIQvL4Cg8vrGtC6Exc0rj6KU/crMG9JAWDsX8guf0+faeR7CreZDyk4RBKU5Ra
Ry5dEjYgfa6JX2unv3JWLNa1Q9g94YuXn642oVA2ud4QfpOcUaw2zJor0DKs85N2Og5BxVjRlNUG
SA199lSy38tljbX7k5TuMWxIuaOR8MLjjfMa4FS9eOPWoVWoK+SMngrrkJn3YzymJ/PBDgNSuinA
+zVcf1P1VQOJ7vyM0p/I6zxSBH8NXFiZYU4dmfm9jqShCatVsy3mKI52EC4Zpj2NaIaToTADAjXT
GJ9iaNqdJgfdtc74pJzJKceYB5zm5+iE+H6X87dhF0A73va27+VN8+8SVwU9fkpYiWkby5bESqlg
KsIuKdhvyHEo0OVOruTFZnodM/gImgitwsZHQmsdN8R4U7YIJABn19dynaKqvETj5ywfotjdXeJU
ND5kJCd10JFL5GBz2SElKnwYW5f8aOIDsmp7BvStBhiyIxQuUfHkX97IxN4qfCxuCKcNKG4F0YXI
A0IDYBdZWgrm35ujRQAno2QX9QwNBHFdoYu6zjwTEOSSgSD0d/NrQBwasEsAnLFzRVrCWqv3+HLK
EXdRF7tu2VwEnBSpDoSAN3dX+kaQW06jnwhA9oWBecKY1OmHZdCGKsPnyZmbqQLDypGXgop6zOwo
xKSRUKWDOtakUrV+VXfV2Z30CdeOXydqyS5peAXbhqrZHjBn/544YWSUzHq4IvvgAmB1DnDvujRc
3UrWz0K4DB/W7dfSpcoY7OBNF3yTKDCQoOvKje5bs4PP4YFCSULZu1Wf5UjtOEa5SkSYJOrEDH46
hnqL50HfzE4xbATIU9kC3TNBvGSMOAb6A4HMugxtx8cCLpFIL3Bmp864NWb4rNjAiyrVaSt60gYC
AXKsjhV6hl1pmWacPWOsQcLV0TIg4pbDoyTVFwDUdCzTBXjhCnBkHmQTuO47vCbXJ3tkhdh6r4TS
74plTa7pXikIPZ5E8o60Wn3qTGOL2EjfBBZzsa4BW7BM7FSQjWF5LPl9FrvO+yMMfbcbhHNCU6Tg
2RQckqC0ZV0jUYHfeYOR04O7+2E9PQp5KgfZN9UARzVHVQfDmOb4Z+xPH+gh+hDbBGR3Tk0G5sEX
NrZmiWVFMzSqXUZsPY5c6n+QgO65/4BSggvsmocFZJ5sJht/BtqWvjsFnKVfhA4b7p3V2jJE65c7
pfHjo803nyQfV5/sE//YTJV8WvTLNEN4hlkXPx5jthihhqxQgOCCXuk08kIzuUYsHp2eMAHR+lu8
pszjZsHW7THQ9A2T8IUJui6+6NiPGlZNM7l90wnJodC/Qfsh8JksREkhVmaS8u4sSfmIRubDXXgT
9Wx72fpfPMT6Co0hO7QYGoakJrt5JJaawKdLTPIrv5zO1oOaLmmlNKNPGXJQXvpSkl0om0qu03rz
OYN+dwyagKoXj1LL6xtiVJR0al/1cZsJq3jr75HT+0cSzUOK2zH9P6eOZUfE6gqCZ0DFUt38v0sX
c5e2/JNex2RFk87mgY2ao6yHJARUMf4p9v5E1Kzzf8m8OYCGM9PxowXd1KTJEYCBhcyRSx5Ky0ji
oHF12fJqNmDlpRvUn6eZ6rOolRyT1qblQZhs3MEDkU+WgGCPcBx85ujsSeJ1p6gC1qkfcfrzIOgV
kRLTKMON+lOPe9DMWfDhxHWmp7ESNG6gh9fyLeNZuMjKxQxxyv9NyDA8lM4EntlDx2y8gRIJpfla
Jhm1EreZSulF5LBR+c4BJa4UKWcGY2x4gs3QL6XZre+I6KURe4LTykvP2mCt5EZPAJiMRev8MQ23
aKnl55sEMq5OXqrCYj+ZL4fz2oJcp3O/bKSoyiNUFfY3QwrgcvJVsk/8I2Yhoir+MIOX1AaCS3AD
L4PtlrYQYJsdGsPGEtv6AQQH7ek9TvjV3LhE4MECGtJdRrq8Birj3VY6sGTlri4DYdkXmd2FZQMo
OWpmsoXTBz93jrGtpicqA34YMyrVHBMdXIL72xAmo8ueg8Iu7vA8nEvt6F6VksTklHIOW6sCjXdi
d5zvu5G1ZnpyCk/6MCbkLHqDLWQhKEyNywJgyPzev5abI7V0B+uPijPoQUA7CYZHM5VMuTBe3Pnn
7YiAHurai1biOc8SAaMFcX+wbzexH/ZMcD5d5IlFHYGT4GhrIHeajC8fk5C2+QGXdNSiByX2MBZA
28STlQ5XG/V3HbofhhincZOEx4kbYUynf7M8rhT2dCQr3i0In8HAsaQ77F6BK77DugAWqkSFxlhA
gc1uvdPGfQQW8hj9c62PEZogPD24+NNqdmyYB+LkatGn8+UUrmt69/eTNerH5J7Xy/OAWczTH6gz
2O952lKPlm9GbATJGKNAEgDrUjsIqJf8e8ayvIFVI9hXDdnMCJhXECH2deZteJnKtIux0WPRsmY0
fHTzds8BLBbBDJa27ZZwtFZfVNtotNFMkTMq5M4Al0XQW3DVA7DuraGu3e8FC+6rrQo8d96TamHg
iPMpeA7nPAqKmP/XwT/SavEGIdRQ9UGvg5JhDeJJvGt8BbMq17BN8EC5sLrF7hBZe4qFzx6jpZjt
j6fWNxanBBrjQIIv2i7xW+2SRj2fJ+cG9jwNLmdgGopl6YiuRQUQay1fKpm5czd2fc5leSqBQgjt
hcniIG4W/aND/SPeI+YsslXfUt8Mn8XPIgFRQobwFERwKgO56XOvQmJJ9tyVCt0fW5jqkvGEfsix
0AYgbSrQzaRezNQiD/427bcsa3sD7Jl5etMrqIR7RcGpZS+deLqx0m5H0EFADuVWLALcOqaIBCvW
oTiXrL7EVFEcrf8pWQW2sIFhFcUlDxBYZIetfIM4Cyx+STiBuwKGDSIxnX6gKcb7vux3JIFs6db9
eFUQzxnkngxN1jdkwIVNT1V1VFWVr0E7+w0RGL3e5/nFkQcwTDU5t2QFhD3+F1FTYDYcI82XvOBM
kE0lXwN8r+f5SRlz5EPIEvcMAqHux74lwFgMJ6taeeQkbpBam0UBjfFiFHW42vl0q4cW/qTF3mvy
zKzcGAWIZMagmc6ybmHFzWL/Nh3XY5yUR01/irH8I9w6OOFCwRAze0VIbVpbJylPYIti+evDR/i1
zsO1YcLMFWCYZKwkCwD1ahuAj5DvP8QWox672DuwaRTpbWHf0gHSvWyXaU3VCvpCsS9876S7yW/G
eXWm3JmjXVPboP0nPmmQpvHJa0fRtbH7UCQ2FMC1noRWidT3hQ20lZzh9myha5ybCCJqdy9BQylG
6j+ZqPSlqr7UWOE9orTtw5fkYMXUUSget97dopyccGbCjBRPBAuSRVOvuYRB67jH+t94zjZB5HFg
OvDKK6BDDtHJfdRQj3LOdzNNPaZGG/WeTf9nNyz7B5VrkYUxksue2URPPiW0d7ZY9KkpfXUe2Zv1
OZuQLw+x6dOgYaJl3r36T5cSclbt4Jm5V0GPoTxSsDz56wl0xMWD4v3bwOcVQZkO137reZ1L5CZ/
ZHpv4uZ2Dlb7fk/yWBDAhlLcQg+/XKMywlklUZuwDdYiEYGW+2aNi0kqdPvHqu1nmZRwDKKk2+4o
BMsWbTZo9Jo8u0VKpic6LVBHAMbdYetnmbUV4X3xwQx+mKYmUQ6dlFJVaUlGFLOHr8w90Zla5NqT
dmVQ5jyb7g4ppLBGltxGtq+L5fririJlcZA0yY7ZA9ThqvoFPNlMPxpZIBX5ZdZuwjYsEmOgsoyI
jGobTRRsVSjFpqpS+w5bTwKEkToMbdF5ER6CfehFqti8k6PsMZqMK4iQvlTKgjckyLfLymdtIjoK
iwZfMk/3yvX/NhwCLFiWaETTeO3aGnft9UQK2OKlNCVhPckKT1xWHDy4V/nE/GLfhrrI8wR4rNxR
JyX5CJ2FV2063OwO4pXUlks0Th+JVKL4DeX7r5dILmK3DHRqwa+NsdGAcJ/wLBRQcZRqKObe7Sla
DKf5feBx7aRrVThvjZGo18ViMY4m8JKiwi3knbSgV0VZ4WQXmqHweoybpuwMDxwE91mRqhuGGehj
7NUMO+mYH9amfXa96TCnm7K0T9tYr7u7tPi6eVt7Bm6np54RMS3jrda5BU9Vj2gBP/AQ/4y2OhkQ
joN6a1FktYWxP1KLgEAeGDlleIUYEw27ea6VUxLwzgqhzjmm7XCo8KMv37qGZ+OLH+L+cYPD8gV5
r9IzPqT4AKIsIzRprOOLOjbsNBZ07N6qpkMnZRnx+/wfsxz6cYP+9nitPygdWNlfJln/ElBAGnKX
5l1T6fOLhk9DsgHNzHrwY0iQGCSJaGXnZJZYs5bMI6CeNdHW1iBhKgaHuhVTiXwX9j95NB8rEjs9
yR0n7umr3ytf4IBp4ZfLnbNvTlUgu9dkz8v5Xj4eZv0l0uwwda2NTmUv9/R1EESMCeBrqUpGCOxM
zEaPs4LKsmZunec8jHYNrAy8jfzAmZhsqD51xzNy7X6HTs61nf6/lhTfbh1fmQdssCtnwWVc6NkJ
IL6pkO2D4jBsrwsj8GQhnzVGm7x+1D/hUVlasAPqvn+FlCCGXpFyjUnHpV2qeYnpvcCT7TpFkpJD
nc0dbLlxbPX4kPmpdw7r0Ogmjy6rgREz9y5nmbuyC+XSoOpcN0O0PcmKTIVh5/G36xnTkg2iaCmE
7UKvDQinV4R7ryamnLar5U074avKeaw5ffIoh3P6z0+/KTAYwL2td65aJ0P8QqgM1k6va9VLDAwv
izeG9lNptoS2wQt0S+kHyk8AYNFT96u+AFg+7Mr6ngkIdi7+MORHTqkA5j7K8BchDm4PeuWik8Rv
CN6yYMKEVbf4aJ6KK4vnb1HLRUigdNEgdG02s9LSdx4JaegDQ7WLzJCU6SZTV/utkAOrD5UBlI25
1JzGCYD+VYlGaWCzbpp7Ud1XIQj00Sqvkk5mlreQnLD4r/AVff90ai+OyrAGY13/2fxaCKgAXTUd
EGIASp6wn2OVGn0+DUVFitqDzM9YKHh/OxPBva1HAMXcrE2qqapzE01Hexv37saiJJE1qtGe096o
ccSbxHt27CXeu6Q0BllvkS+KEnHcgBWLuUYql7FPfuTTWsFlBVbbR+whHGs1IoZ16w0Qc3cqXPNO
RGHI7ZNFVy+kT9frF5JDeI943hhuUhaL9w1A+bc6/IgJAEZXgV8T8yTyNDMMWb2ti+nBWZh52hWN
40UjLC5jhtehC8F0MVSCONX6xR+6SwYKyx7A1Pjuh5xP254oHzDM0wzKNDLlbrr3Fv4j10cN1qPQ
nNgwQ3aBHTblTmtIbn+4pSSBNimxQkoB1P08Imr8odDpgoqX9qZiPyQFjjGyNbsgaY2tMF4wZZBc
i5Tn9/lTAuS0LHL6xu+8rbHJFLGU0d907NzZ7m/mABoVLRMC6n/p+sP5Z3geEkfkixbMx2tsfklw
cXieEVmacc/YOkTq0whFS/cjlKE3SL+RYsLjcXjRcFaApzDURe6dv7eYtxvQErf/cNLrP26yxg1Y
ttWR0IMlqUbvZGKNWvSWHxrCVatKJdJhF/YNifl9NLYvWJLsNvF7/Qpna1zu8Ucq6fWhXjOvLmNU
wqQo5bJBr12BB2YGFboZnSGeoRPtDuyuBeMv/FqcXDOuAGLe0JCGZ/SoU0/yHp6iev9AidBycIFI
NorhWMKG3KJ760yWR30xrmyc72R7+vIeZPOpvx9kFZL4UCuc8qSWQZTXhFfUToAC9TfxPkJmZERK
vf17KWau8tyFLstoDQTTBAr+huwWBMfJxxQ7uDKx2dKEWxOeDcLTeE69j7/9HHjQqyMd5RAC5RIW
DXbpUjwigNfRFJTr4fXiT/Rf3ZT3zlDOkCTUltQq9yW4JsGBxLnLPRKG7Zq55SiPPbTl+xLyNwPp
zzEdfkbUe1d14vuQ5UUkSPxTL6WiLyhlD+aasRXonTdVzDCJytKDtBx2bPYODF1EOFCz+Bf9FD/C
8dGzOJOqd26LbAQlMAx89J/6OAIF76G5njEMINvJSQVbU+pKHsNh+BYHQN+mX5Gt9h/V+bEu/3gW
O8oVpHG1eQHqQcXRCKkdxL3fXEOG8dnvMp868c+yPFvIv7RlhDFfpFbagcAzbPWQebQDiF+7b7bM
qZ9ALMeEUM2z8G+JyOI0KKkzn42aSsKTIq2l4BZn+FDiy5zbpaS0EkROFA3ohU9BNMw/253ZcmZ5
vYfoB1/UVxl90Kwi+vk3PbhLH5Zktbn0W+xXzYAjb4eGmHk+h0Chx18xllNsqiGC8dRSEMJq+dqT
6FmBLZVO5SHqnLFZu/2WYQ45UVRX/BgIvVVLkaSUx+cHqNeMLJvbvQvHsy5uYoFcF9iqTWfEI2qs
JqYcVLrrw60bFSO7Z/yZCYqPBHyNppBn+p7cc0P5XKrins+PhxSgvYMx71fwbkITwHT9vOca0IhY
ozjEcNn3adezIhY3VLPIIdAfLDmj4OwPddBrBMpgq7uxhHwuN+UOD1qTVAl/DwIaUxoBAz4GiyeM
Lhqa22iKlveDuaTNA7cU6gGrmHqSb1W/hOJ5PoNYTpwTRkScTEF0xICvB+4xi9xgEGYvzjGf9DO1
0EgmqBE6lxHRI0PeZjYZKWP3lDGgD2rCkIa2BHUR+1jGLzAWUJRPIPqyA8PGZ7Vdsn3OhYKHkh6k
W7cdkWCex6pGtsllIwZCAGExvf8ma8rhfOF8EgEbi6QkgO0wmEX/XbC97MROjBMkuy4vnPiphFkl
ixleS+NDdIqELHOt8896NYb3k7ecXSE8b50sjhioBIMvOI8WmC5HUudAJ1/fh5Xok/DnhQrW3CdZ
xA7gmczvaFTuDBvw5TTZ2/CXWIAGevk/HRMHJj+iM0D0rHqA1d/KNsT++kclk729ZSayn+knsidI
0I5HWr8AHWd9Wm/mNJUNasF3eo+ERxK6vmshwZRLarZzKfXBjCBhrGeo8BAg8k42b68PpIPqfzlT
H+zBPznuHerwsreIuzhCKAVjXt5sj8mxBsOp346DVfHDu8qbFM4IKdQ55pcuhvK9XFF3vESS4pwx
QPBIfCqVxg2IGXgnK5QA5vHvt+jwpnjRB3UTFg0nXHHRnp1UIxPrYK5QiHR2hWE1HII5/WmWz+w1
Wsw8oLNtXbDIKwnW0pEJaxajcj8fvVZUek1pJY7fDc3j1Olp69HKxxFe3ZR9IANz0RcohW/6bfaG
sSsk46xgZTPRiEdokklOvf88UzD7jNPNIMvtKWxQIagy0HcZ7JFX3+6tFg6vSZyo8I/qkv5G2X0g
hIoKSAawKf0ayRXAkk+/C0A1mkuMm3+58DKJwpv4ckILEpIGk/dGwcVs/sR9LIdR2l2YKhOf0N9w
e8R/xOob4iic0fmuPFofAzErEvAaF0EbkhTVFtYd8OqngoFqUVG7p5P8kqiD2bJWV5rfedv+Qp/y
fe7GFNW/4NqMFywnaJWKbLgqMFUFg0NuuuZh7P+CmNt4YtJG0LQiYeu7AvlQXxadO+LJulpi/ckJ
bK0KPOuF8RSdprHEQMA2172H5+ThoCWrR+qM3zTeqNZO60molh3KvauZN6VGHReZ1+cmpBrRBJq1
5iyTsqiiXDTnnrAGdhF+qFOsdOADdasmckQCAu1qlRR5065UjAGHihXmMVrBXpHubVQGz15S6Ll6
WczS68LZyBtWwvjX8Eqc4vdQbMFHU1fx0YVlvKpAeabc3YHhllOjVj4MgfukMo+fupvkE7XID+gR
PIVorJFzDe9SCikP8abEeUfDLsTrmq61D9EkgOnnyPWvyw5jJTd587uAZZWmyhMcRXjAJA2hglxG
68oPkp4eVRRl9tZ5+HAPi42GwdJBojRuvBesxxYz1pzZsVprLhiHCW4GJjwIuxAzcomDGxZRz3Yz
2BESMgFYo48qMy3qG70Gh9DcwyjeVvt71nkwnni57znesNCmvvvpLGnkXHFJluArNv+1vTGTtPNT
blt71NNwk9o8yWGlc2OTgqkFgjQgzL0iGSTL46Cgk7Osew47wtzoHiJXdlsZ5q7xiNQRgTgtgql9
uM8lzyetTnjz2r+EO3gYxa96ScLc8kwQCUqGXOUVnXqi+6HTJNiN8x1nPfWfR7FA9eeTmtNQSlt5
uxZR4uhSYNe9x3RZaTmXynJ7E+IYtDlTCwuneaqUFaKo/5WOhxs6pmsQ1Ia09uArnzj5I4PDkF1x
h+f4MTePSO21Oqq7G3ThGkZiwFRIoT/tMT8RV4yqmIlHTUoNYY5CwfJPFspaAA2o7iJoj4sxiB6G
Wl/BtZiS7zQ5gAV2DJuLTBUvQTA+Fn/9Tl6FNCBOcFNOTFW2tYHYRWKXNMMhMi+ot17/TbhsDDVn
2JW3dihBiJF42630TXi1EuXRmH6p+TKiyowVcGcDlDVMcX8vcgG5gza3p1Q+WogGSJbO69UCnoYr
uytOsU8lhDxnFB3nvzH6myonYhu3qi+7ScmjIk7qQFJxDPZg8UINR4HyU/4Dy6djel1YAnpqcdwo
hrFiIa7iuTTvG6qj8DRI1LUZPDghUr62jkMWG/eNFjvbUYfSlY0GIJs1ru+g8G0zn/HTYIeF6NNQ
uyGrRJV35v1T839JUxpajfHTVtGdZd3uHh+gIJ/Z9I2axDUn2l3UwmsmfNDEIZgP9N+M8WgG4qZO
FkUSTezzTANq/fUKd3YqOAV4jz+b72V1ZLnA7EY5iOkASMT/r5qb2zhsyGjJQUO8M73UgA9PzAIL
CpekuKLNwPA84zmYKY53qmwD208c1k8svFqhgeVsz6gMr7qrG4bd55rSAoA+vaseqkU/GUjpubaW
/lHIM2rKgZeRJ0gNAgVS36UZrDwpEXi1GcATltERwpTQr98gJqXqw36L4cITGbiyCu/jjk2IuEjA
0yc7mPyNTeq34aOiF+qcdBI6S5wAPHdUUxAHCUMQhQqZgiSLQDWul5JwDFM3vnqKCnKpGbBNhTdI
44l9/NetHMHWzjqIYYRiqa/iOzivJ2dNfw6futIjoO92H6wTZcxhhPlAXc/DGoCRkL8RVeJP7j2T
vC2P0m4ohYIf0NrEu2y0VZcKF4UAPxEoDLvJYm9PSyWNjsWS1WaCwA765N5pqpQWBJO0dZj2lMBE
YB1Hxf9+P66nfdXPvKG7+erDy+6Pe785RRQTzdd0RCvLLzhBJ65ahF8/Ni9OpIAVd7gIwC9I1D1f
7ZO8prHbsz9uwRBbzvHyG4z5PZij3Y3waXGC1wnNwqZom0jgSqwFPjKEOfoudSNkU13/NjhctkgH
XktBWT0c/n3ip28WEXS5iRjki8dH8eT2XO60ySENtfD+MrFPPAr58KlRAmDJHF/50HnerfMBGBHR
DGvekLBxguk/yd/XInZ9d76y12Z4VY0Ym2/A9ayWYaqtusz2TwXc0b46dBl68hgbWpFEk16bf19i
avaH7+sjZT9XLwgWDbWKmqURfNzhfZ7LrMIELlLsauPjZQ72QJ2/mJUEcUr9G4hp/Uvv2mV5tp9U
T8uRQV3Ni0nYAtU4HloXppOKFDHRIttheMOmPBVKFrXdGPfiaoJiEEnb61e0Lf0fSYtA4ADht9zI
cRzXEYO+pVoWSHcNGHOy51ffRuQOKkDb0V40Cbu0p+2A+UUp3+IaPckbvizhvwnyDA50fW+bFuWG
wR4BORUHnKWiEB56qZ5z0NBHAjq3Hi8NnRn1orbP65+0QSeL+vBhO/ewZxSxFCwlZZQsl9NQkKV9
rQNRT3WwPO6JQfM0XmjHCJvzxd6o2ALVY1s2HPHrUYPFoFqz3YHw8NxN77q4o57sGDiU4tLy4zOK
rL1DTyyP9lFynHIOabWktqV0Tm2lJXCqCUMgnYTa0Ni2P7XzPH2micm1vgiD7Hi5Bd07a9xFdF3+
tLu9jhQ0kJaTNjAheFwDHNZbNfXECVsmMIu3BEQMivLwZbRagDiudvfyBejzcZG71TzI4exg0jok
83PjKYYEaBM2x09PatOFK1uqYCaaJkco9Ioq1y9y9/j/UNu6T48F+dPOWnM+tFz7sfXT0zWHdoxT
t9tTEerQbAb/iiIWVPiDIxYZocZiMbgiSTPeWT4+0RjjtoeeEFYIg1iCbMwZu7a8Jb2f0WOnFeu9
bPawnVyfaGXNIUNHYKND5dB5/Eg4scKqY+TmqQGi7NCZxFPQ+bqsePLmD2C2smeob07JisyWJfq9
65tKsDQToBS64Q5lYpdMmtWOW3+2diHwzT/JykPmFPlvFAfC1MSIrXQheZu6z0XjaGjPOI50e27W
BFebnxQCTAFVmQ7HSOpI5AawlWRo4hFeRi9rly1QzHH1+Wwl0QHvhitHDjQ8SFGExAFPbTs5YfgK
/MuAmT/2xAa8LCtrYMBnBN2OGkDtpshBLGxPTL1PZK6DmQvJFatGZkQBBXJgTHK6LY2iBJKw0FJ2
mt1HfatQEwostZrprMmttTWEPQdLWB+qeTnSU7Un5vrwtInbaXRlQhNoTCRfYgAES5o/h0Brv9TS
CIe9ZF1waT/XA6CdBwCq4Z3F+etN5d+sHMqdzOaDxrWaYudI4pEz9HPul5ORqp9kHf/rHTsNEMbb
5OLMp6Nx+3OF2rrwOt1dMsQnkmuTbP5E156Pcvxy5wzEEuq0pKd2Lug6sNn3OP/7b6oX97Gd9j2Z
9C1IagUXBWxf8eDxRHtMaRCz0epLQMfOyyJO9z9T1T5F/n0741TTPrpJClHfr3ymwfgptyK58DLw
1qjTeYdHoPMiRgTzLTPFieXZjKeJ6OFIInJ6lScgnwWprP33AH6zuY0Ph3wL8Y8mJcBgftNtV5hq
srxJgZ5sY1pDerBllWh59/aRWiicUpJZ8LwL16G0TFNmM9phM0d4Y7jIOPFbwHYqvXMkRyPVKEbT
0QtzVa0dWcT3DDli3XNrF+NH/tLVjw45jYKuU8XNgYtfYU/iD1R5lSIUgn2NXsS6E8HzA58Va7qc
YnS8BxQOiT9Hzhd7Za0eu89QRD/tdcAIV0zvO/jaIF1SqO2Mh4bq7F8avlDmoRXHzlTwfiBBsybG
kg11KDngPshY4wYJBjc1WVaShrdngb15fZaBqX9lQcPaTtw/D5t/eD4vxzxcTc9gkJzaddH8gDBg
8HcVd/7yd4TW23w4icH4GHI2gDxCmF+u5GpqK+ThJ5bvTR8cV9l2Xs8/tz7CmdmMXwDk/GN3mVav
c0ZD89FqecnqYTxydWM0bAXDWwhLyJ9cLDFMckLSTuFP0Tj/kLj2a282A0ZF+GWMzJ7aMRgrplEW
3lr6lkggI6GkOQI8pFceQatV+7MZHor/NpvGX2BnTnoCNKjVsyad7BilF8NjwwMqbaHFnxq94pS5
C0RzUbmXEGg2VA7FkCyy0pSHZMne9UYXFOMaptXGIrQ+nd7hqbGqYdPH03K7+RQpiLd0octCUULR
sUiOPtiMO28rB1oI8vN5l0u6gzpT7MjDp+SO2P+DKYxAbmG0n/NSZ+lxDu1fVtXZ7ovuI1ThqEdI
2+jbNKKR20BfDB6H4ilz5TcPQiv5/GB/4J/mnUzIXGTyCGBaqos2GoS01VNJBsnds2adoKEBieoB
/otm5Ztfo9H2uCFlFnnt0iFbMj9+QPn0Lj20/IYw/2Ykx1PeTc2o9Q+f7s/CAOSil4g77dCyq07D
CDKL2itqmCGipxL/n0J5mEK3CMWQTffhMTJYSpgp3qMzvvdXEVn8v99XxemSZ9kvcJ33i4ymas6K
/VKnb+K84blyaRBidFcz4DxcEdGDt5yhjuf6ARx588K21ulm3EhA/jRpCBlnVt8/7AbqEl7O1zjg
8ZVAThwYG9d5XtGJ2Vnl4tsUjtyx9CV8MafReaP6warhq7+Ds7hhLUomQhiFBtOdcfCYczGE7Ggv
m6OOcOGRJvz7cAzi5w1bpdB/mlkTgGjgERHLbyDCnmWuiWmDN0b5piDe8S1n+p0TkL2daRHAPcYU
F5ockxCm9z+X1VaVUswnfK8Wgz19M3JvmLm6ioFTTwBB9n5ilA3TVQ+E9C4DlUwYknc80yH1uhOE
1u7xlYGWRGmfXQOq73lOjW6ant2BNDig/EsrwMBfSU5LJKIJi0bYHsdEpOwqOIztAjCfuInxUNnA
p9eqePZqzgUny1EEe9bdkdeiL0I7YadRKVJGN5N7nVxaW/wxmdkh66nUKnkLBP7m8tx6SQ1Ntr7P
fBr76qC+hQS4UJPWGo2QCsj0UTDzfctHFoUSY93yCgrBvElt9Nc9+706qkkHdihlYjtsjzVH7wzT
igjRWiK97Mq5bd+jyzAUcRWhKwv+k2dFV+9YyEqHhv5O76EVUl7H3DeZTllrW+ThjklqMw3xQ+oA
AfXlUKbBJM5LvTX4gwngSd1FdZ7oDHqFOpSRvJTV/r2BzoFl4VN7pU2igSnsX2lBCk+yQlLQa/66
jko168zTN7f4RQAKf8Wxj+C1GWL5vq/g3K/XY7BoMNz2/zxVCzVm7fuusOdQSYb3m3Ze1sx3dmU3
km4Hke7tOc/xTaYqYhon2W7Pl8WRF+28nsRyVhun0Uzm1k6UHLvhNxffAD8bLKl3wkc8crek9d4F
a6rNzWg/uiflhdPJFxiMlrcJAsoD3cSvwZqQ8YKdOjqq5LZ2wIsp1RVjBsVkR6F7yGXDiTmUeJPm
BMy97nhxamDuvMkKz1IPzizrM8/ZcFX0CL/n0b7j9fDDZHTDhkb0Tpx5H5oqpn18v4eIz1mGMm+D
EFvAZelWZvBRr8CrpbhvXtVvHSHUvnqluBJ0RT5d/MXcaRlYSMJOfX9T5VVA1WgyoHDNVMu0ja1V
ofrxSpQ+kF2i9DaKegKdlBhJN4JnlDQKjllWx56WEYWe0ppd+UaAU/zJ9HjxklQ3Ex1iO6+1q71F
GBi0vBzsenP2MQ5/DaoTuF2s4EO2MGkfBNfDPC3pkaxXcGyknbgyTUy841YtZZxjRcI6jWwT/E9U
2/9gzcoQBLb6Y7X8eSYugdOqbuXmv9d9UlEL4UeYmZqDdTCqw/drQbrhD5a2ZCYnCliBrV9+dSSp
38xh+Z9co4GtkpJ9MtwO52bzwDEf5fC1fsYKv+G3jPzH+yHK+ms0Mqte85g5ybLBhp1W7cFu8+S3
2SPF7zWU/aY1qNtgw0iCMOSr8MwCu/rQadOhxY+jgpuT1dauy0R8u8x+SWZG7LUSmvUyopxO04Sj
RKAah2Dw0QoV6N2f5srSbHk+Qztn/ChixjZ6RFabwQXPd1FF/UJf/0kRWhAzJYewaDnggadoACBd
hzVtnV+IE8lHdjdCF4kHjuwrOvPB34lAKIQtelvm1Z3Xo8cOnghslPUrKBiltzBcuUtzUyoGAxfb
fLuM8XeXUI2R27geNNYbNK0NCcm0wn8qhMjeBmpxi2Qk8iQ21qja65AzZvgTxywWafLZ8uRzggHa
Jiaw83mg5K86Mp1F+M/wWVzLhMu76fd8JZmN4/WN9wHayYQVzoWlJb2T8T74kI4G1IzGcalArBy6
xh3O+O+JEuuEY8lhJ/qObOMVa84iptEAZMiwYukEoBhYH/6UGi6VBB0nyO2YxzzKRwtmFnmMifL/
1HXiH43d/B5wKH2IWpB8OANemPv/XQCslUdJgh6fCuxahZVxxW+DHrROgaOeKm3qqct+q+moW//8
7a6JeSF/RQW4YE6jN3Yr1225avldeozAEwd+UUVVu+B5/3BaFBwKK6D+6t4AB0gAQrNVks+DcSpa
gxvbvVDfrFp4yhwH1ofyG6J7Lpvuh5W9HQD5wQZOBc+dxjR/MHzvgwd6m2zry/BaY+9kGBF8hkAM
W2+Sx4xVAxuTwIgC/Q31NGIx/baJNUkaTYTlgU3XAxwS55FcX9km9n42UBqefBJAK4ttY3v3MEOq
TjPWXUFQl8dUXAju2kvyTkwxkhHKNu1D9HtTRvZn/xXGwMwG1aLQScBYYwxurPwUBfHBgaw8GwS8
xexW5nPsOuTg3YvmOAQ/++IXTQUETvy/zBs10Xk3ol3TVIMUutk0liSxlwGiJ9/qhEm5pOmhV4pw
mU2LyppkVeRPFzzUw59VyGnn1WIgsjBrm0omEMH/q212HmC8TT8Jjalf5sWjanm8SLBx1Ixb7P+m
5D/li1UyJfXrAKYDIvx6bTQtGSpuy1Aq7/Sd8mHPc+bzSIQpRwdwpnomsGzeuBDGZ050kNj3HK+q
rkym5jYhTkYYRNjXr6mVsDP2OSW9xkMKWKTAcGorzXdP25/vPkVJY2TvurzaXK4nzVBjje5OplM3
PE4gJJvnLzrF8nalbUTB3N1mRHfoFOKJMT1BlZMpEhVO6dxCDZSdRIgpaiXHhog+higg8zAOJ2Cy
TySDi2h/rTOPQ1Uwa8Trr5mvl0I2zenwFRgOweQYpd1BYiw4qG99e3qVgpaq/bHDF5KC/cr/SF0h
rD+Uo90MW/Vm3CZTrr6bC4+Si+i5QrrsMNCxSNJDLxnDIOjCH/t1w+UnLqnv3+fwgyH7QZoS4OJ4
r1WP3P27nnrXCn2hLwnSCYWC9gV+JuZtMLOy4cNNWp+rN7g+l7vahNuNJshZbLgUD955uppeA3Iq
EOB7mwNU0N3abFXBrMxs6ccVLrzdNUTk5yaQCzgl32E6oLvm04N6MajBsNrXVnXx/4UvC7zSISGw
FmRxePmREPQXnmQYfCZozLW9wI4PgGsNszXWe+D7B6MRVbHiwDk/2Qw9BCn1Mc1WlRJpuhA4Abhs
3ySIAAd9AVFNPm1q/gDUjY/47jSbcmIeQtEGDWWxwHm/6nqrvHDHh5C6DmKk6WQ7gWyRMxy7K6Qf
wYsdTdC5KmCr64Dp8mZj6Oy+8qXE+XkEGrQNVhe12jCp9Xyh/t4Wb4/iv6+gpRbqBcWaffjQXKFw
3M0WTg8fYoFrkpPooJTzqHLvX+JkBZXKSwjIkSN5v71+UuxQjogQlGntEpgUu4d99qwrVd19xXl0
HChEshyPjY6YCwrCNFjTzoJ/chxWnY51gXkEqQpli7thUqtHzautVFRL1j2bdaPkX5HbYQFUQFuP
s8i1mwxEHjVi91YLTJtr424Be2CR2IJxyJmKnhC4Kn4sL88T1ve8U+XT0D32lulomQmEbYh9YkfJ
z8nUQipow3jurMaQNiNHPD9/IdThtrbVszww2OqMlY11+BDNoIyKAFuFVmljeKnIyiLeso/1214S
QHfDbNtI4sSCAq/4r3ML7a8EQpuT2tgm7tSlWtoC9GtzdBz/lvvCTBQ81z/9j57on89DoL2tBAk1
n2ynaT1I7n0+6ZK6iwzJ0R5l4XZkf31aWAJY3NhyAXP0tbPrJP00jLBRnAa4sFTX1e1mP5nUxKZB
Re8NSrYP1fOFhRERLimSrWeFEqxLZUcZUzlhvV50I83XIRgbTDEugUO1gg4XrrUVr+ZdRzlzKmAz
OwWjCs4uEnB0lqcxqRE3JRaAZGZL1swqRpycYU5H2770fwS6zC/8cLlO2Nn/rgklegEpLoDAvi4Z
h3e3UOkDuAobSI1cBqe6UV1ZscGk8M/tgKONijOtUSRNk87NHJcsTGN/gDaoSA9kFthDIM4lMWaJ
lvbvYPGHNGdM34G+kHm2QW8ga/kFA057d7ojj7a59uAA/4aY6ult/BUPSfyaG/A4IJOGVRWuKdgo
K3a4WQWNzY09x6yBDIOUeqQWWPn9mpvgE7wDKW8VbJg86Z+oAMJljkKYNS8uWyUitijN87goAfga
7IcjuBp0Yg2SsQqg3FoNEj0K8P2gf86rV5or4YuUAFloFdbiielsjTon9ig4dG3ZRZWxdfOiU175
c2dHKBovkubCq347/YAqAEBRVFPlEae/Ght9Q6DsxF5eP+9PUYERxDt8SltxX43mkRqj0oT6fIhS
8yNcQg1P4itqZd7HXAMPSpF2KmhHfAPTLAf5K1CC70tOSZY/K95BpbHZXP7go4TtZn/4Mu1lWyYu
naBWV874iDjjLI/H5in2bDTTpsFYIwubfhLxGnfarVFs0PUrnIWmr35SW/tvOwhIXMQOLhOjg0JP
AWmeeCMqyqFO/TA3z5UwqOyw+SxC8mqz/fkhGpLLfWFF5xdZBufJVf+MUqa6QBydPMArF5CdDWim
QuqU71d11AfPmCxjrGu03I3B0FmujPpiFxPsSBbJPhorrz1uJBdAdL7SRQJxiLjXdbD+cEl9jYbm
ZwDPk7AmGmcqWRKINUZhqctsZiOja5bipOv2rRGAEVK1Wy4DBNluKcpHqQDwBMMdhN7D9yH1UjaN
tkGXchmqx2vWd3XWdOX4L2e9KhqntS1rVnfr2hFxQgITkB29wYZIlnTXbw/YVGUBpHu0UeGC8uw/
mVt8R3XRmo8GrhM46twXaLr9hpY/ATFdVKuCiYnCkOncOfh+5mNz9rKos+mLq3p3cqvqmqgsE1X1
s1gyldt92NzJn3gzpaNVGegOa8Sz6e94Znz7akqYGLvDP4QTMyJiD/3vxqQ7gEQvpEDkxa4qE9Yj
FEUkejf7fXiqrpy+FEr4LegQlCBhX8mbU60MT/AQFs7bq25E9ScSWBI7PdAQVHdvfFBHMBkeZpY0
mVtJ7N/UHT3myjwjPlq9GA7/7nmMBAm+7aFXmmBJ6LQXHsBSUxEvgg7nr7lgJMcpfX/W6lofCfh1
aMjP+grE/QHSIw6PLI46eJ5zLKC3Z3jCkc7OWZNwcaYaf48GgALlplYvI1eV+2xUhYtdmdVzxyXG
nq4IfFPXFfYE3Tmi7MYCsmhd0vxkPb/V//cDrtmfzwa+JF1EHcYDbAk4+w1xJLxojgbb8k3Dwm9l
P0j1Qk6l1VzKJdBYkcWg4slPdmgvkuFGQ2WGX4hYsHxIwQqQtR66GbVF2oYJMfcz0XNdI9qlFjac
IwJK/VU2dYqxeP0YjG6fAAMN8eWktUgX/zCNgZ8d/yYdD/FeKrJm5W2BhwQpJgqO/2oEy08FHB/z
rcuTpsc16C/ZK6tdqDGUsMQRstmRaRPJwTXO3FnZlzW0I7VJsSOhNnmHAxYLMQ06CHH3whGRP+tp
/H4i6TmyiX98zBYiNG+JgoVcejSlBUpz1idkRD0gLdzp0RRjtmcz0Uld6uD8GfjOpq9udp7Wd4Gb
pWATwZcDiEwv55nGstRHxT/QT2pKWcs4z/DcJhD0xJaw7OmCHEMm+EAcjaY6EyBmUKZg/HZtzZIz
O0dyylX3cSS0T0gGhktpF6eVJwKJgTGyD9f+q15wHyrI/LLN6CgQ43ZxLoG2zYCVz75s9uwj/K6t
fpbpOdVFJC8BRLtI9CFXbnsUYdPp8HGnNlKTakoV334SmmEhV4js0pBI7H2n6mYzByzD/F9jYa7E
3Gl/Tnv5oUwYDmozCdq5GP/Rv9SaHlsf96PFlCKHU2OZ/3BzETo4Ncj6sVih+v96IYyQVal3CUQH
ow49AIx/+gFGS9hcFwtkJaxFehy5VjsDNEMTxIgOgr4dFhzhUNKlaLTxub7pqa5DLjZQl4XHpX52
YyjYhevRlP9iSnW9fxVv64Aq17/O5dVnFNjOJCTcJuDfM9z6ybliTXJJ8mBVYD8/IwBTBXhO5Sej
lRLL7EH1F+a/Eh2ljKXJriQdWB/2E3HETYtJDRd2p2LIB+4k35XFDabqELpbT6JDp+a6F86DEcOB
jTcuRwId0VeStQg/4KxZqI2yhq+3wMfAmxtPyQvYpXirtDcZ4Kmhlh758A933lN0nZjtpzZl/w/v
O4t6U21pxQKL9Wk/w0nR7WKI8u/gX+xC/5l2+fPld9K+yCcLAq/4Oy7XXAM7vDyX1Ecmvrh8JQVc
S3ZPGLK1IMeorBakO1f24dQnwfEMwqrNvzVQqdivI83ShGNxn1nbU4ZFg7fkvlpGOVUV6eTZv6Y9
IdNeqhGWqs4cwvJijwEvXmFrAZYDax8t4+kAnQIm9//O92lhE2NuMksZomEu5EW3L4UM8vFbJ3R7
yktQSB33EVchnVi76QCJAkpQ19WPRMsleVupug9XhtxVLklFoSNoI8GucXGnwRS7QLqAL8kO8mT5
rrbP337xhU61PpkIeNUb2qXUeDCykqE0M7nkA4Hro8FCO9v6Df8hRtlxFEkdVa5PQtXih6t5pVzb
BdW9ijyhPQbU2mqdenoBD+1f2so3nrBIM1xOj2COP083XUy3DFkjPJ9BbIk7PLYXug1ajr8W/yPJ
UEa0Y3wI88+zRDx+dPOdQjC8LrMzrNOSVl47S4k1pGStjqTdGBKRDEL6UOvSwC9MZdh8oQUlmK/K
J08OmwSicipXvzYplQAfXypkUZp0eMeeK6M6OUK7FnWcpJndN2aR7Ocf21L2HC3X5RbWfh75wZht
BFWZCZVXvA4ZtNZjS9LSpJog+g72JEaXpw71/mp3PDvVwUYzfm5Uo+XurH7qk5VjOBz8N+cttCc2
jXMAGOiLsjssUzw7MOsgmKNVist/s8F4bc957MmM5NwIEpDSukn3LFLDHnhOtJiyfqCAq732ep71
+44rs5et3X2aGBCj48WhW7EMRWYEtctzIQ5pn9OvSK8ipSbt8+JC/AkRoUkXDZ1ps7RYFzQ8fkTT
PUcoasv/uUJ2lr0rsrj7B2pNZj+0LwALhPki2KvcrK+LuXI3330xB/HK57dmsPnxTJ9CJzQSurQv
phL5Nppmr1G2WoHZ86zEd7JMXDPgD9d6bdQYN6Y0vsJ7tBn7viLNcmc6mxAONapcTruW3jGnQmkB
XgEyZ4RlOb4g/PZyeMgfy8BlCwb3R3Xc2EEMszxRKNOy3tM3DEU/znQd9/j4XiBY72iiaXnBzHSQ
u8FNMY17vtxbEhVvsq+oacUVPA50ZF6THatgFSejXGOEF2CAlNY9U8ZfXlDRXKZWSlMsPYoTFzpQ
Fa66Yctik3iy9CK6Nc4i/dIR5uYe30nb0l+RSxnsmRIt6lHTgOUMyYk/Dab+Wh8lyePSzkFQYMAj
jj0ODXVewNGOS0K8bkq4UdI0Nsh5RBtlPdCDUN9cifIvFIXd7nOtcZAK6xeugxqJwEYXeQeHubhk
XHAdvl/DC+wL8JyOJT1Gayd0gSaPVJqYjkpGDrEELjDFGgiCwi45UVq2QiDDRJEDrT2Ksae/iKxG
pucUKOHB3uJSG8qCXJAx7EnJVsoPccDIl77HSsZFTbO6ky0RY47UvdoYoJacS+kiLFNVy8HWw8HV
4IL9INrp9/VxvTttGl5p0wSATwX7VXERNm2x14cmng4DYGg/9+pNLOz4wEuXPuVeriuuOX/Cjznw
tcPSYyjJDKXdvZMIXvGX17wUBifFwu/Po3LVCHKMrR9E9bDIo+bInAsrlNBHm3NUtFgQGSGj5aUK
8KjjypqktvHBEVkcbIUirytDYOZvAud/Icrxr+cccy2PN9Pd7iD2GwvXvsagSC8Q7grrFb9L5TMg
pODgHj6zOmLkMk+eDsqifRifCL4p4haTC+u4AkIJRw14Ezmxwkfdh4Exdvrsgo/4ArXxLHbwDyvz
csuJ6uC7V7kxukTI+Swc38KL0PfAUFDJsea0/R118Hp8wonah4vjc85g3MtiRtz3IwBnYZVw4okD
REwg/cduM1LeEZcoU01Ds+euFZSDI85H6ekNJM+N35redYWsdCVOHYoZXX2jIP+U8kDjS8VJt7en
ltaQ/5XHzc8/kFcKI2I1JfJCRcYuXmGu1K691tGq2uZe0OHR+fitTbolOt3N5hZZOHs4NZNj3rgA
+Yd7h+oNYDTMZNwYKZCyPjFmfwqJTrslfjzpz24ubMKg7my5JTIiyhCO3T35BHgcvM83DiC5Ap3j
20DjyFTQBJCUU0Ys09VNgaHbFoy9O1D3KkrXHJTv1+Ezw/HVVFvq/eqIlAT7qNa6w9t1VMgbD/sj
ZcLbK9eBFf1iA72M2D6Lvq4iPtKef6aovkFQJ2dmTtRuf0dLG8FYdyZ3Gbq0XnLrKgCVywKsoG0V
JYmcKRD8df6yEzcRemLDaRcuwzLSULIYOAf1dgxQQj/z+KU8N+H86NkK6GTrC4koa6URH8eKLKOl
lGmMeZpXkNcLEjujK8Utca+q9y5qU56ZeK0OxunxAlBvJfJMlvbkER1+wTEbPbnXj7PyeFsOVOHC
A+fMPMDCFz/2URlzPO32ziMkMbyq4gMj0JNFcft4SK+7GP2J62ZrTF1NRAsO1lfR2FJ8stEaXKVz
BPK1buDMnFgdP3uFaf7RTp4A0YaRhsJxTsUrldx71wiB53rTqLPSt/Z7IcJjhxoDGQsxVH68/u8Z
rSpz1lM6fz5vlEZYQmreBjKeGcwu8CWv/fS+rNIntoDumNQOmaAA20J5Z7YfXK8qw4anAKJCXxB1
1TKEMYu3BR0X0fhdWMDinpLNpzAEiZrY2bWS1AiBlq5WJ5YaHqe1mGS8k3Nxd5vGOqXEs2SfBzgL
VJtJ+P42ZP5IkBs/5/taTOIId5koJGBsgRIpz/mQZmnv67l/SJHCfB2Xr57dSLa9762s2uotM1Ho
AznUngDviGX4jIIEWh4i8RTHs0ZZbqmmvV/tFt+7pwzvrDfsqGRNskVNWBuuSjDjSmPE5f1oqZiu
1vaufFZruB559ePl161UdAB4SI3YqHulMVfXJ5UHPfPuHewBQhlUqCKUM0u/L8pVar1LO3quxfP6
nECkjMNZgDhsrfcSCegCNQimN2JWrZZE4MvKCFJOuDwxoB/0L+Qo+MEcQzRXbtOS6S7qedDjafBV
tcSqkIyNtnZhaEBQojamzjrowznsVOPRxLxDJqEsUBRPcG4u85aFTadKAo6rQZYU+nm/pA+XDuk3
FvYQRmpnG4ocafDBIyCD4mgtIxsHTMY9dVa0cEFtSZXDBXJ1+G8EHAerivHWi9B81ZAjHcObtOC/
c+4i0GE5rjc9SO4ACmPpG73/4DUkdg0F3SXC0l0a2l7FWhYKGUGeZ36FRZFKsZr4aMhu3HOEYqrA
kOXgUqPZg+Ewy23En2dE6f+a9zXKJv7tB2/j/N6tWpikZedXH5NOxCwbWmg/Z01mKrrtRKjexwQi
kc9IKrNcftBRaVAwj7xgITcsIZOYL6X5Q6nf1BUc7mOoYsjZCOyY2ZiLMUFdglqmmOTWvpt1NHXe
EU0WdTqJi5bDvUNg7gDCxXBcgqkR0mkI7D8uMc1Hwv4SoIZs5zWsrMIB3KuN5MDhMdxTwn7NWLxS
yKyVP/uyOvY6aeL4a9+VVKnERk/CvwfHOs5FW8Mc33OFXg/mq94rDWXh2jP+WlJNZq1qhD8aKhAN
LoFHRPQw6LZ/MPoEY3TfbSpW1W7tAZRuuXPMqzGqYTm1jWa/JTHIu7JMA3aEPn7iybzDH2YMILDB
jIsFNoZYRnA0muXX12miFd4vzfhnLSVqViM8zys1ejpC0JxEmzedZtSTseN5KYSrpjZtZ2IhTnQO
aNJi7xf1x2Gb08ZhbJKId/tCt67AvNMxcYE5yl4XlxscpQnw00K2DaYBEV499Wxpo9rxmsDwplpt
ts4MztLLwVuWAcCw0HxW0koje4o9ewhnyg45No9FGsj7npLW0aqwylqlZ6OhTdbk3mSHKK7+ltZA
fJ4Jo08lNYVFvf/rGjGZIGcZ9wMFV6iA8Q88IAv6odz3ySgW4HIdaoLKpdflzuAoBph8f42D6qzk
Fv/H86BDBeDzj2YnJo4nbYbdXJWBl+9U6QgSrm9Oo2vu70TX8ao0bkdepRwRrLRjjIxptBbOHsNe
UsoqrjyW+FdBwQ5NZfyk4dNDuO+fPiMZoZr4JNZ9U8/fF1qwUOgM97Yyuqc4j7q1OArZVhkdNuQJ
dMLO0qJ/jCdjXWg44rTb06hAA6OFj84LhtabtwyMS7MP42x8hzjsWBAjR7jkNaHp9nX3qJXk3Ipk
cFk1kn0Jju07Qq5UDEO6G6qwbuWJ+ifB6ozKg5bk5VUi3os6b803rJJ5Rv3suixe1d4eoLj5bt8M
dJhh3RbY5tRs1WBghGGJwHA+w8xEFHbLXvOxEQO9dB8z31sQKE2OKkv7VJFvjXiViTkiOyF0Mj2g
6Clk13E5lh07uLwskwFARwWCnmZwjLD1yV5oNWZLTHOw9nnSX2p3lDhqo9vOt0zr0pe6u3394HoW
k1/zpKKlZ25gwRVali5fcVFjlPvmdgKEUeYsjvfHNIVBwkC1HbolpU6RClrf5OcPMpe5Q3IF02mS
EtZtojRsB/LJrDaAswMAuGImzqjobjJBqA/OBJ5n7iHnxHuzYl3Bg+t7kgpkXb7cYoIAosaMWcNQ
UpILyO2bNrIai2LmZddH0cQwmXzcu+JVR4jVsA0OW6h/tgovR2B7HMgaZZyS8OZoXBVkKmDLZOOZ
DX8qGem7B82fljRxP2EZ3IXK9rx/k0smAg2ChOYsrKv38qlE+jIgVTfhZTR6y5wLl5j0oPOVM01L
975xiEZiTPWAFT6rTTU2i95UMiWLuUoqW9bQm91i/3yb2rFnwN/bFDl+zt3x3UQ/eyvhU4RQWWT5
+WL7M+Urz+w5RHJOZMLw+QSHZRrZWvkynSANEFFO0F8wNCkIhlEhypa174zyHrWXAio0bTLKTPEx
LkFCARoQ2z7EqSktAAhXhkb4XaGNhaAZPiDvcXg+3iW6Sjz334+8bMXJWgyoV/2MoF+xmrdq2Egx
iAp9YYJz0iSo/r1arbgNSEHpiHeiJQ40S4lmeG06ZcTRWh5Y9DhAUqqiW172BowtzHMI7HBWy+Pf
XetDGfD2f45NaAC/zd4+5ogEYYFMv0G5PoWIDG+fIRpp4qUS0x0vSKwHvPy+ldqj0Z4yhW7ZSxuv
oCT3PMIIkkM061KSOkhT19ThixBBDw3guMQ5gq3iEI88sujShhJrviXF0DeqVz9PjuuIqf8mFJYn
9eGA1Re68mQlOw0I+V/ErmFHydz1Ka1VDJ00qcVj8H1vB15Z7j3dwApFbmE13Ef1xmuy0NTbe40o
3xrTA1ZXH9TGEeJ9yLzDTukFPmJXylenZZUDddH7+J4qEUF7oDaPWTsTdhmoFZMe5hZaVI7wadm2
rPiSJju3FlPHC0EyX00rDE90XUYZN0zFFq2W8o2y7UAG+sqgT1GV+RhJqCpEK/90v1J7rO90SJae
OaV4DWq+s20vqV903qJ8JXbNLuAv0uRoX/ro/9ORWKnQhzopSavHaSDkOorY/V6oWUXL5L2kDYaj
6OR1xx5hQ5oblWQvI69+JPzi3ryLnPAotiL0nwLW/t6u30/L5xEJ7rF4C8Uq59ytrMDnBfCJIDcG
BxMwAeqcnDyKnCx7e3j4+dDGe/vNkZfUMI8WqsiimTxB8g+ps1PTwU0+wL9OJnmiJ+hQfzTzfNKf
0MX1lgC5YBAOCEVNBpC8epXZ5v6zeOx8bxgsGYQPHMJ+5xjM8fEVgUl2et2ypK8EhDC7xi+MlXnI
pI+X+W1Hwlz2S0nNKzPyUdV3c5TKRcRC47GK1h36OOXfHl8LdMdSlUy3zPswZedEAHmNtOXE5exK
P9KHiT09AA3ofppoj2IXLmGq+V07wHbRk7KUDMfkU89jlTvTbrrBEAiN3QrwwYoZcMa3b+m2BE9u
3wGR4w6zxQ2UaJ3cWcZhnEK0oCoGPC1yNAuW55MQiYfhyhk3HkWUQ6QlZPYoxY7MMvrrJ21lOzgk
i5jYu3RK/ekp+itkJmKtkfsgb2/67JYOyDpxv/4I+0N9w92E2er9cH9F9bOJUGYMa7EHkL0FDl4D
Nmny9ubHrNSCx+mQcigyh7+4doNnNvFvWMKITkkJLSWcr0P0LcRO8lGZazy0sF/3K882wVH41Pml
++rWvDMWEIR0xskqC9XRWMG02oB9osEOFLM15WaaMmNqkvnvV1f6kSJ7+kf1DoLO732sTRC08DCw
1unU/six9SuG4feZ2un1+VSNity/qnm3SLR3kZOwYzIO/4ovyCm3Md1cMXXDz6baxjknVhEv2Wlb
3hDYuSFjsOmNqL3xb5/sFTw9KylCSnahGo601L9sGJYuarWDBOuXKXpL8GYviBHQiv5j5fyNTusZ
v/30B9rwdooSqczXEzZgG+Jxt0MFelJJ2/MfTw9Ng3n+OypdjYS1zHLkPX0q8y9oFaa/MuoEU7HV
17EnSxJ6sngdgRqHmA/O9hJXIo9KnJ7HSluBq4jMO7U1CTPzCyaNQLwmfmxWmeHAclfy0R+mMO9n
0rM1MlytsegjpOKUczHx1soNXQ0NRqVGSpeBfGsQx+GmplCd5cweVaRtwBXzR5tn08AukMtjoSSF
0y/Sz2ZfIIQ1dO4avIexmzOoRaVnMnaEu0mxDMncxGeaqMcYJagRDiCAXBMV+HUVS8h+pfovm6hv
Y7aDf/U8/vLjurIo4RaJ7ABFCDwIWGvKziHMD0tO8vrvumHn7cBtd4E8dtTgPYN12oxL70NlpFUV
Re+pKdG/Lh1D3Ig/TcjO/fez6Le9DTeQgqSPAddoBNsRAd1mop6emJuIueTf96TOQIN0YtLDtgTX
pZOxzKCvpBFLj6jENZlM5g8muSQKhj3TREeriCns0Y+F1e1NIaeRmnzgIh/KTAV+jF54+E2bTa4/
TV68SKtB/w7vGM2D+JoS2ZyvfZl5+OMyQtg+qAJrDAI/unjGMwA3fjdzKjw5k/WptHyX5LbPXztJ
BmCpmSwHR7RyZusPRv9/difgaQP4XAYZJMXY/tXHH2ntOIDKqKNfsYf4/vD39LUgSOYWauh1B+BQ
BE2hnYl4+XDpHLEWeEVGyRsNQRYuFkDO2PB6NT2dExbyU9D1xokXrp1GiXtjKr1hKQiEymnH8+9j
rOTIVahfoX2UssW3Nnlarz3/8pDA+q2oPEVkOANs0+3P7jvno4qmyfZz+k02dOhLN+wpV7FdC89x
3EelV5HFGKTflwWBzMR8hJzL0ONObaGdbGztnS2v4RqRqhu3fEHHEu8mgxrvO9fZUJR5s54wP4Cw
Ge+aavScAsV0//6rOsYtoA22YjadFvm+N1DQJvIgtqD5dpLmOQbo4Fi6qQT2S3KrhyBjnYZWLZ6p
tIGUpn+ue2obUWBIdOtGJpyGeUpRj0umVg+T15c+FAI7lqpnZMmLHd6sGNlraqPWLbVcmC53Hg6G
tZq8eS+J/gEGkkIZm5zT2SQf298kwulX3DzQc506t9zlnNWkxZWhh9/FN9ZHzZF5JmsInzmy9hC9
8SH/eCqRV2thM29l46Rmngopa4AY+QBu6WUad6Ey9GVE2A3I3yxE5uQoylH8Tk+lyn0U5ENgCA8Z
QZMIPDZ2uUFd8JU1YnDDUzPbZCbre4MRCQ8kdcn1ojm1a1vaonuCvKSkLp4cAl2+liM4Zkqu6Zd1
B1NT31fgOh04+hGweeqg8Yscu0G3DmhqjcZYFf0Bla4UQ8PavCjdn36Z3nCqgfKpfaHHl/orr1FT
tguG7NNsGJd8f3mScJKp1Tzk+Y575JmqxaZCn+ZCaOwbbXwB4bu6SnHhhQVrbluEEjJtOqnqdrYW
sIxHpLO2ZqdV+7+4cJc8BTi39KKNr2AQXMA6PWJoX8k2iaDaERGi0a0ERq+fuYAaTOuU1hDV8w02
8AHjy+ZCHQJ45HzReTJbX6Mvuu2IesArWN0HHJtl2ilAqttT4y7rNlDyL1V6licokNVZhpWnbvel
ac0U16tLd8MgA8y3jKc3iC/HVnc6RwKMtbmGMo41mqLfGjnbFURgd5L3Szdc26OFjpSZU3UqYaIn
xXCzpc9M8ZUsYqosres6+ga8qxl3JFOSLjALpffiCD4nFNUXXWZFiqQ0bzsrlynvJrIW3BOhSZ0k
aR/7RZPPM4Utf1DrCZdrskDg8W89wYmQBsNudnm59ahLiv0NUYNl7UhwYddJcKOzXq4VUwUTr1fd
iRZf3iY6fjftt8k0IyVnPT2WFPDqV19NMAiTPbEUcGEplL+fbStLcO/2xhVPnoIuZkuxXO+L2HaZ
E9QeANDr2neRCqNrBjkSCx/3+uzttUGX6/dN95bRcBoSVIU4JU4OCBgEScazD13b8voOCb5Uj7gN
D//FOIBqZF6W4skTy9l4Hsh/MJ36Cw4yJiN+kNI+zgwb8MBz1/owohRTYsu/vEjY7yuqcjc0Wa85
CbyDqdDYFzn4z0joxxIeUiGztympN17I4Gd7rt8vmzLEtfyf8i+lKSi6dmvrT49ehP7q7ay+VuRm
24TSrCtylZUuA3u0HsR86tqu19uwH3HQcSqdX8ftjPD/eN+23rtNXTQEfohbMifkJF3qR0P0Ynq6
2HYdNAeHl59iqmy3OhEom0EDb9WRavx8KzGnVetnffcgK9TGggMTC8BtgeUQ4+ClOHHLqMk90NqO
iCPUNamoZjMRO8J2+sLnJVinwfrRZKYz2997H3IYyGIS/gCbEpLVhEmuYbNIwGrdZUlmkl/BtiGa
NLLEI4NgIKiOBfuUxPjnQLy0pSMtf0bE7twowretRtWWc8aYSbTFVMbXZJsjlleBrjyQORfjhOZC
amzcywBVEisGq5B/uoYQA8SPt2SCzl20k9OMfe/t/fzSPZj3DxCLQPms3rSod3Pzrp05mX6pXjyP
bt23fwFSmMov9oenaYSoVOgbv9b4+8bJuyENCuT62Oj3Y3N3DMJYq8Vsq+iAEaJd+B6iV0XtQ20E
l7PkoOR9xwBGA2AHlbeVVRWb/aHbfG5ZvCyH9kdqoEiYRBXzB/X3m/ekX24ZfOwlz9ARRklYXcL+
KvQsWBxv4Y7uHIyqR36NnglVra/Zhr++wDLXDMY3cHbqq2z6IHgxueR4R4B+sv1HxftcgMd7Nh4b
irPS389Cc9VBp901Tp9Ho/sNywDUl399Ib9UlxGRt5QwWzV+tdCBAdZidqgHrdkxFnSu6F8WxIuz
VoCQKjopUngDA8OhNzGCuTayvzK1tDvIpj8kt2YGU1RLvVURxlFr8Ir2XSy/uRS2bdatB5Ul8f00
fzb3HJPm95srw2HosQvzuzAQ4zotknVHfx7w1GY5x+Kk4HPd3rKPyKRcetwekYsd9u1srCMIvFXh
OUa5s5bRT4ex8w8NPm6UhcXEXHx7+0miZYmTpLTH5dDn13Rfh1Xu0WyCbwjGNxPPNfJamme9+imj
fWdVEPFl4cTlUg26Ema+Fp4m/sAHbVBsby9ehPVn1jN1fw49QG6BI8SWkvgR/Q566r5o3jKRWS4u
gCByYEkPkWNxvS2df/iOtfA5adIHGhgQLGT2zflaMthB3GWl8vlR92EUt0kTeHmfaR+QPByWElef
FW0Q0LTALoRSqmr+Dvf0AmFWQvJvYr0LQWX/g+fPb1PExeQGvGMm8uW3+cka2rlW+HEZOrfwTH+V
OjwgeqC0/VZGfy2JqxFQ8pOzamDy8aDRxI2FJF+3K+G8+hN43htbZVfCluIT0X/enQzgqpEfffqG
ksGnS4FurZcufZpHMGBt26Bvx0/r5y59XYTBTJjIAm+9eSvrzVpzQjJJi4mugQI2kSgqED9jhKQZ
oH5pjoHprMo7Tm1CufzvUrAFVdeVq4/r8KbahDVQRCXEopmBNv1CtB95GdvoAAx1xNytwvUzdsLe
yn4dZqR/NtNTVAt4RVnOmjsTPD2KAiW0fjliE6YA7qjc6EivKg8wOmwd3q2PMDHMMA7gJ+JnWcdE
6vOX7q7l8No3AaNc2HU4xchIrZlvs4l7Jw7dO8Lx99kp8IWjeZa+mFe8u1kjllyIYh7swh2Jmdua
EEd3xL5Oh6auaaVKdi8qb/eVfSEIUj9BBMKfPF5rbdMN9Af/nAXQ10bt7nXrSZ1//cTH/HUsiK0H
fqp3Xj0NTRnqYACsPHjArNHAS0aGlNXJBqS0Wvd6L8ZIBhAz8nLNRPPjZf0vzxpNgP6pfBGX8ynS
WHHyuklxDpMjRJvyxrYwpp16S3+2YkOExj34Mwo49mmMZsoHDKfzd+Bm026gazSdMNfVE8v53LCR
cTp2Y3GR6cBfQ7Sf3p8cu/6Yiauba0QRZu90FZnzUb3w1gEjePL8HCFMGuEb2NuVBJgSGS3/bm97
HoRbljD4If/ChgfwXM6LsM2/P3Qj08sc5/pPwGs+aVQfOqjYemaehWhekfTue8Hd2Rbdk9+QhMja
/vyWIM5SZGSIA4KmaUw5BbZYmoMRIbR75MHFVmhf4N/93uos/amgl+/+/eiVMx2vdFq7me+P/qVN
UwkORu3CPuu3V6V1fOUkYpcHTq8zp+jUmd3RVimK6wzVPu4NvlfCyJ0JbAKWccSB0K6T1butp42f
c7aAjel0czEsP7+2MIijj2tEJrgj8q4QgTiLQyEIx2T8bwahALEZ9MNuy8RbgFu6IdG6SB3RWdUB
g9SWwalEkCguapM8Hm1SmyP+gOxkvn47N0wllFdQeUFxIz3l60O8rsP3lYgzQ4UJcFT0XHwm+AAh
zH/fEQq8g8ktdYaf+xU7D4ntNYO8tGNmZmYcK8FmVfgNCC8AexHScFbvFx4bqDeCYeSkkcmyQQg9
AZQ+iWShimXeuaIF+3sXTk1DJ3jTLZ2sjoCmgrlYgRxsZxwFLFbkpr2p2L4TspMG+t+7rSuZ2w8Z
CWGG9VYQUAQk6IzgQBmDozV+msk4zvGseg8ARujNlf4cySOtfseMeTDUHEsZeyrKuTqKHpnLQ/RN
HHCbW5yH8ekSAw9KbeKKD9Clp8ZYT4dJd+K04PwgVkrSICS8iHsNxln0FaoT4gH9N/PwAaFozkX+
2U+ukYOURS6TfPkj55+tpq1kKmKmWR8TXxR1ANrItVttPrvoDcB2K/mQ+cY6Horndg+T7tFjk12L
AyhrZQMHnvc4DjN3NWC01uVHTeOKD6QJdP8vpNqePclngOU3U6URrKTX4KJmnNVRqpY3ZP54mPcK
6Q6/uwS+1RRReOelVIgGs/vmktFUCFRvxP1Qa5gs3+MklQpGYR5oZpj1rMnGmsvySUR1vExKrdhk
LMKqL/fqOHBXKPhKvtoQcEhYqzO+cnA6ApEeI0CSEACysWBY6LGVh+ado9CJiE+awjRc8e744mM5
1uhVInpP2B71CmWbOCWyqJNZrBNFAf/Zfj60k1OkKhx+ALp0wMBrp3+NTc1uau+6JyHCppWttKS/
hnMssvp4RwuGI1mtqyJ9C7DH3fC1IjtrPoAQvigoN+i986nJiCC6Tt9aV7d8e7N/0BbQPSmbK/MA
T0uVfjQUU8IRHx7x0uLaTJjP6q3Ya67w3kpfeuDQVtLx2jPqIKLxTI0vlR/ZQJIHXgtomByCoF5H
awqJNUCjTFyNpZgl1vSzMu1+p9yMDoHxWhQI3rxrx/goqXMzoc/HK3LVWTIztg/2llhH77pI5h+q
ajjWTp++3put+Nl8ygXM7dXx+FeNkDFwsAef6bG0SLicP4ICI/fs8hnl13c5Jv/9QSPaHgYshCAi
U8wtVsfpu0QsjIKWBJZ1ezRYAtMWH/g/zbk1Dkz+VribzZMUA/lK1nyglJuPBL08fqNY6v96LUbg
3jli4umCevMbWtfUgM1e7v9T95PdghvDOWB18CsFdYURJA1ixlTU2SQA4GLALTZqVqRT/2ts9iCg
x5uCx189bttlH2H7IOS/CPJsyYjzI66XaDZAgQAs1LRpIDJD+sa4KleFZblHjYEnHc9a96I41yAE
KdoTDNSEJ0pkTEo9qoCwwqk4MoPAPyC4ZHJ7schAPYMqt18D9JD2840FZEk/0YZR45KFmPciBzrW
m+slFlsnGc6P4cQU4IV1DgKfZ+l6zUJxo4g83mZrxa6v1gC7AlhwCYdrGKmq25LKBAP+73Sbcn+D
kkK8VVmC3TyT7hV4RTJ2ziqJmvC8SDyzS/Tn3/xp7OQVFzFR2lmeS9GzvKugBBfAXAVQ1XacP+WL
OeaN55rgLJocO0EJEehaPY3FUSU+nUtlhXMoGKFPASWtd7z1MviSppChPWQZUKCCRXK1sOzwzRjN
hk4Nv2KhuFYPskIGlC1zt0Bl1THHHnJaOhiSv3eMOS4YdEuhy0FjmUQOEgUvTeHR914O+GO0hOi8
/WK6p1Tnsq3OyvKXJh6qnp+KtUmqK/4Z42onjZsfe1JShcVTErz86AuTwL7+IJF4z8ByyF+9rrRk
R2zRytSNPi2Yd5H7a5IC7/Nk5NrViO0p6SHRjjD2u5wd03lpVZ6A1LaK47fnUmMPLVmC+NxbbkZP
oqPrjFuhMosYILPcGb7GN3AQUW6GTZ9A/kltTKmWBzzsO7fj+nyIPpyh7VlxiMU+vSgXq5WfpmgF
jfsJyZ1QhVyKn6ZDUDvamKzpflY/hJaXP4bJftyMe4y48YxnYieI9KKB16iNHUAkbMPiRlxOtR5W
uBHFtaTUNm17AANzThr/qITdxFKwIiKn5lkL4hck0Z7EnSU7SYBZPR2q5aL/q15dbL2qMrK1/HzN
sccrruVeNCyNNIrGOR6vZjGfgtLL3Oj0Y6FGCepvk6LyAhP6dC+4A1LLf3X2yQ9lba3WWON4IhBP
7bwSLtNdlJ8trSNh2P6lBeyANLxtmBOwiuOBnDK3Lz71NbL0CbCTTKqPCQq+Bo7Af/fSP844x7Cc
bLakMskS6lGJd1uKkFqgxOksGZ5bM94yH8RfcwkfVLZHgsPOQzzPRt6WdKS7FUa0pX59dq0r2lTo
eobRsSrhLkzTaBo+FgaEsT3r2CBLJCLSy+ENRMdCyrMWMgkYF+WywS57h2TP/lgzPKIN0wWA7v4V
t3eLXK7Mj95YEf1NVcdz4kT0gtkGseg83B44AutVK0ZozwjXaaCHL6i7HfTwdiqWv4YxrpJTc8Pu
f2XARj3EQvWWXkPhlt8ge8pWX0+plyymiIz5cdQacQu/teZz/xgDu6S88O1RjTEDQuUnSwxPSBa8
fTeCzDnrHtBxIiNVQogJbQWajO/zMAFOiX8ih8UYtvWCyKIoewW8Nu1FEksIitdFIwf9oUYgEjUo
bb+Rv61u2sqYi/b0SZytST3iklL4/hxz8JRpQM+lsZsxX8xWQJRVpdTeyjALmHpTezgwE6EGJHBK
fxEr5x0uPCmHevMKZu1H4OnTG6hj+LQCrMnDGjXzV4GUwx43qJoIb6wHVuJl+p2TppqPjjFVkFMq
sNabTydjjxlnQ56K8A3xmI5W5XYMsvx96WqYS3QDUccOdyDfmuZoeToMpg9I2g39ZipOrvQyrfMm
pX22WNxSoKdYEBYhNE0LPI+4G6FA8XYztAuDg2o5jWMr3myDbqx3UboWgHDrgQTqLJ6oQQoudQOL
uOyn7m7oGH/u+t06KTKs9cSys6I05ydRHBieAzd8UdWtE24ZECAtitRLPUWZxdnWdpeT2Lb+u1kX
HD9UmpBjPaM/CYLYqmrUSVifY5wwymQBqWhUQwu8eOmso4/SsYjo+SJkd/igxbIIx9XRtOF2wJJS
vUnEhiCB5Niv/blPx4ERvnj1MNzWQHULTzrwXVSg+qlZPQIlpmgeCBr/NfCyfnUhcv2oJs6dRKOr
rMh1zKugl+5mWf9ejdtFkyCcpC6prkJxByXkmwIO0tiWMGjoROnjLMbrJ45maBplR3tjj2BJ52Sz
bUApSAMSoE/uJDmXMdPtfA1I7L47tAv8QknzvYLnS5fFYeDRc+KTujPcq8NZczkIko1dHWN1+oi/
gBpNFTuQPYA9I3+8oIPRD/iKGc0+0/9yy4LfrfU0Yfgvv5UxIV8WcwZFCVSb9uAXtnT4aV0NIlny
dOxxMnxpOuytk9HwMMUGeftIxwXPZbf+MDoT64xBf/eAD18fXTTqkL/72t5odxURaDbj60w7RA7h
DZZ82NufDwImmROScNlG3W7QF1J43kW4GUtkWDriuW6XRpGQdpfJk8NABQDiSpK48dh2ZgquuFJB
eLIWnslD06l8/mnJa2TXu2hptskSUbrzYvv6vVJGLBgwLYs4wIAfa7+K9C+H65MmWlENIFkwDDef
m0ZXf9DWLVu7o8G8I2WzNiXnZdlbysbWd6FZTBYBs2f3+e4bSjlrIc3befnEwZ2zy5xVK4GsGX3J
Q7+4H675ZL3+hjFDkRYuyAzKWlptKR8BtHftD2uKt5GZtDZAnRWnN8nCkr/Ep7c0O3BBWT/tKkqR
/RLGu9FZYU8dEzmvNkl/9/w62n0eEmhK87KTpbpB+cNotEUGlX+OWyv74yDNClTVhErLNyxY7Gr7
y5bxAP/o/uWwGL4sf1wp49713/Ndc/uWMEiBQnr0Fhv/Ji8ervZBwrKPvDI48XbJk7QM/mQKmCgC
8VpE7WVAt7g48z7rYilFpUbB1nhO0wtiHhRAST4IYd10NWHd4XiCtP1D7wPiFO3xJW3ZIajMgisG
ks67VYVXwKmetKpmW8/XtDjGoBcG1Nx/Q2T1RWzhh31oF4KjHRVjoEXk0AgKO42EKJOJTvmtsa70
smUhYEYzw8WfiVsxqcMSoHiZd648Ij612TbEnsMn4lfmI3hz3Gp0kI8aLUSW2RNVHRP4/ifgXqp0
+PAcpeDQKiIj3bdnGOqCyoR6Erk1JGKSUREEiaHGBOdp+I8rIRjG/wpjdMEI0k6+r5sJLOC+1p8j
Mv4cgwnCgLqAtR7GEB0QTohlqL+Ola6WXaZgMAzerMuYREp0fioMNrSTxOepuk6KZzsIqMGKghbF
CSWg0KAkZGl4JqBqZzutQVS99cBF9QZclv7RDOhsoWI/Yb9oLh+h/nUM56mVC/2UaRy4a5LVlyK6
TR7cz8wTUiF81h7+2x7wuA/SB30VgvRAdfXZI/fKfmyf+KWuQrFHHw69CYkYdbwfdySq+oVd1BfV
z6uuXLc7fwQ/50DEuk19+c5BMp9jN/PpkFlhTOV0tYBxTypDpdvJKqBdY4C99H2dZ4RGkpZx/9LZ
juR2DTTH3MGdTDwNLFe9xkSjYlTrjmmd4L75sErQtYmAA++SqNalvkAgKo6Fod89jbNeOquLkzqO
Vz2PT02j7LDEPP5m+oMvphQGwOVHgBi5YMLeFZisC4RA+w2l+gp0q63gQTH8LEaNQ5QeAE33q+GI
MnsMMJKXjA1tmj9nwEj7RzDeI0gl7qmcgr6GdrsqA27oYSLVXiewqIeZirw4BCol/h7Zr8+SvSen
VYYdLtgCppcoIhOPrh99lrjSR/iCaFHAL1PqNIGFCO1hpSq1r7JBHVe24gaaq5XYDnAGz2Y3alNy
KgXzh7Bu1HD2iphe+x2b00b054fN+/BnpplLRmwrmG3kOMRddVpNpwMBAq7FEDRIqRYHRfERmuzb
XU1kpTEgPCUVUVnf9Fvv195slyS2o/diwpH1x8hAc2UFciyg+ZFiQSvO1AHjbO/i4sj6Plas1lwF
jiF/YyXUuhWGtZ7wXwwSNTUI3M5Nl9M9f9tXYb3VZCYnhgxprk/WDhQh42GqOCE8rXtC8G8R2cyD
BYQ5E9BTaqmDhYe8bFmd7oFsvkdRqMmRTRKymJh4d3qwLctEgCKFsjZ+tpHMqtSkpUc9v1kO/eCA
OtEbg6a14TuVYyLtqKkHa+1Vk3QReEELMfVMpSvWWeV8EyTqZe0/MyW4hihM7FBWEgVW8u3anhOF
eQYhA4U9jGBR21XVisufB55entqgvklgb8Gqlq3sVH/sTlL9AZgTJCSOfU+0APd+Ubp4+Cipnt0v
fFm0HYZ8ti4nikBDtuRSr2sU23e0YC22Ss6zDHSxNu8Zhd3LJ0bvx/qGMR8JxjCE11E77N4bBP13
SmGdOt0lTcxC2q+GusziYjAcENSLvLZDeilDgP1l9/vriPQzVGgCRigjmPgdOwAFoJ3VRWga6I5X
Xt3uArWULp3f/YRvcJudOuaSpFNCXPZRMtWh6nX5iAugTR20wVfLDd1zwTiRQqC7E0ZGZPke8T+/
v533gptyPDbSTpI7ERtaihT471LOQP2Q5HhtedxZlOFiyGrrUWG3DALNMYD/TnoTNlEEPHwW4vDC
q5YyNKR8xPbBmievpfZ4fLqmSntIQ42RVFn77OX4sVKzXdND16vZ7WLRRCdbkK0WGBweZ4bZvUDw
JPcwQetduph0ko93ve3SFHNSDuCBnkshqFMnpB+KvpwuuGmUX3Oyk8VKvK5snKAjETQprPtrUlws
k9bRMnJp39aK2ZEwRISZNaT3fehrnqd8GdagDLHgwk9DsJLA0E36AHViXAFxoUp1AasfueUeXod+
GV1cXBFQ2gzTXudaYewVLDa78f+JKorsAvOTKGkrZi09l1Ma2J2a4S2WNX/wVZJbwTm3CDFq9KBv
ipALFn2U/ZmHqj6X3wsMsxHi45QYme05EQt/gTszhxiL2a43i9xA6uRP9zySl69ezIA3+Ecgquh9
EhfkrUIuhvRRTq4p7dZWO6EBZESed2GOjOkjNYte85MGNt8b6fr6uGcCc13MIhs+u+bnEHALF6Zd
QL8DHJXnqSnpmErlDtbGtKSVjKlrpBOxmL6kwaW15PdlhrDFVv+ILDKEJc17ta3zC8/zHaPIGt0d
vhSxQVvjWxAj8gFCNZEk9NtB3BTE6z7fRmDtHqbZSEIly3HmCX/0f20gbrJqgSXuCr+YYvFT3XWW
LyLbzZowhzuTBLkPUBdBAHlCHjSUiaFuElejNvnwHHLqZ85SeVE5fNS7kmlxRnyN7sMR8IBYm+98
jW2y3YC0OCm/Zml1e0u53KuRrxvpUhOe9RZVQq8XTwZvA8JHkYYhoonA5XnjiuazR+a747cZOD5p
sE1SVxBek6LxyG1ssz4PHXV9jAr3gTmY/yQn8UBuj4Tvvtn/DlHf7h+SzqGGVxtbXp05RaWJKnQp
ysRxKz89Br4Z2BRbSFxfMSB+tM9Wlg3Y28paU+jhzzoWApPuPrcjKhFgsa6aiE/1dcmrfaMeFWzS
sakCDFxTKSwLAvYAtz4hvVTNvrY/OUHiXrTEQxs40Z7EeOe8jx012xWJMbPogJ2HXTNnR5XAM3fc
qtMWTFtIaR+viUQ+kMm/yRi4b8Fgz0FxjhblqteU/zsKrNVM7ibn83GXG02Xt8WAYAZAUdRZ4c2P
BeSU76rNbaTa35hXerWZj7yYef2vnnuHoNnDYFoRXk45+pN6ttOCpHiOhtb1W1JJkqwuGS4Bui9h
zjSrZeU/k3B1XihyK8F/ceZXp0yoc23BlqQFmD0RiBad97QKPdL+LSziVdtF9fAETuYno2lRSjHh
Or3ZW8KU0AEy4rKCJshjqj1OUYkSJ2P5krlQ2she3saya3SA6e9aYk2+u9e+0HDkVlEenluhkFIg
izB443EQ3X6eZ5u0UGshKUMvUvloVrCmWXfLPc86ua2eNSbISIo5zgzmHWOaGyQphED0bMnq90f/
3UvyXGuf562AXuscSspNDJqBurqIGeEwmn2hzmp2okbJlJuEXKN+aMQcIavIopdX1at1QIJ99Q9r
gMOQadmzOwQCSLifLguRly2f1ZITTN0cbBkTM11mF8cM7eovvOZgzWlrLFr55kVQFVbNT0KTARtD
OdwquS5YKsn0Fx7Fd/YvfNozIBWmYS7jJco/zWXBnsvQ2bl1hArWIdH/Ys2mXyXNS95G7XiQrGzF
89E2sb1snPCLYSvfnsFXjzy+Hhb2WtsalqovKKeljrNiMjpzn5+pq3T3g6YuF5RRHJlEfP0lXXnq
9o79JqKkh8Wbq81m8YCytTbTUQ1cq1AfxoXN6Hn1Ct/NpjouDxj7uJ8THL/tfXvIlyvD3eskJIng
90ljnlfKGeAcXNf+0H2JdpQ0oBc88wMVN7ZdkvA0rNNNbzGDu28zALzVoAKbvll0U7VXSi0XM5O4
VhsLO1oatMpPPHCHRjl0BdmdmDBOrOEA5IzMwte22nHWI3NpGXsHFtwXUhjXZsfkroPUAvHh/uYZ
LfvyDd9Mxxn7LEmGrEmeXNvS1La+TlHPR7Z7Ygf8uspTjVYAvKup9UyBItaTcoRLM3aAidenRYWx
MOj+wwxeeSMBvdZCzCYvAVQc+Zp/XwsfVvYxt5TkxUC6W2uCn1XwAHDzoeWx/g8FH1TOeeJ0MIpl
JHtsbRitP657RuY/iHotppbpxKCCbOi9dTfbLQ/wSCaW27+Bpq9IG/xpZ8jcEvPodO3jO3WS18ei
DjXCoPXEzAFjiqcrHsNaSaSIspulDNlrkOwp1ZniALdBSabgE89CpCe1WnwHPds9wYRzEzE4+azb
/9vSCGHAi5EP1EzlmKbCZaaXrzRK1+EeabA4No2+JCq+cdEkZqp4/FXlcZxubegc2zCC2cAFqVUa
d9RJ3jCVmN+VDzn70S00uQhJL5B/t+06TAf4rwMlfVW0lS+9oqTCYTxEI/m6HFsxHTzEqgV5m4cV
E9oVBgxp2PHaI7EHCQIJBwaCPfWXBdM15WTNBhGNH5XbU0hRoaG62jIAfrn/B3zwBKVgvWrVBw/8
8V3N5bNBRDmIH6HukOWpGbI9spNr/gJjl01YOMNTW/aqEwRrhUad3VtcSJPkLvfsrbcjn8An0AYx
AuPjQzdNgk5/Sdv01mGNu7I6a28HV9ZfLwuTNrmMcb63qocpxUpEnOvStb+S9AGNABwjM/QfuY6N
QQaMQ5DVXiywmnjQCEhrzaKQuJ+Ud0mD7c6bX+EjPNmvQxB1eQ3453DPu6AGtOLz372vWuOnZs0n
EY3/ckHV98Bw57Iq29LP3EoI+IdrdXIV0scddfCVu4NSsJNu7KdKJZ+JmjnK0HCtzGCf3VeFTSK6
yFUK7+VZedC+ED0U/9/p3sYoZ75bcPnge25NDGT/KSGwY/22XyZiAzDdOdC4P8ZmBXEuYY3uO1CF
tQ3w2131FN1wlOqzXC0ivT5HeYws3acMNka3sCypdPBuqu9so8jNe697z69mv7ttEpkdAOftIXV5
80BfF2awvU8GltL1UJru0DJzi1+sADM8vGRrPRPf8sC5j7Wph9uQQXaEZS65dGqL3xuSg/7uesli
VRZWw7HUCiFS+W/wucITmKzZGEh6gTR8Qi7TfGOLSuuyJWLH1iRibNN8ggYAPE1c97hXE8tuo8vj
8jFuaEo8wNapDW/Z+8ixg08NQlNZ39JvLCO3HgZt7BKykkR4l4gk7+3yJCeHDQLaoMPI/wPWhNiR
tmEa+K9D62OqsalW6ShaFvRojHi9HrXh9GbK0sLM9MFG9E4lJiuLktZ74SlYPcwey+C7kKujqt93
GzXxR8L+orXokXP8zAUiTxNI4aJKr8kiXlm9FGfSgL8x4DnGOV5wPLV+j3fLU0rZsZnGY8MGmen4
/PGoSn0i9RxUpPNoaBbCyDYvbTlYGL6q6SnbSmNGLHejuYvCL13h8tu41MKMuT2F1S0HKSZGdc2D
ubCgOnhHsxiXPoGUPd/qikOBNuDGaE8FJ+QJsrtzIp8GlNPYKNmBDgSDfTYbm/AUoc27UZhjulKG
MtQsBlklKQ4Wxb3IQX8zyybIqbPfWZO0XiuP95D/le+JI6FFalJDUtS73egqLSWi7iYz2XN9y3k/
xR9WsMRcMZW86nForqwm5YnRlHSXURBD1Sj9CvLnH/wzbgkkjLUwN9FRVRUYnZg1l9khcVFxbeXz
R6lXvSoZl9r8DWPDvVG+ai/0EsBPblHcqupLntvbS4SB4Wk8vBVNnCPPor6KQJM8u3geEkjOvEFP
ZFZpDT2em8DP+rpnQy0JPsSmGnq2ehxzAd4qTDBjEtHEmJX+yfAr0mXdbbyDv/ihHr7EqXpwXs4L
J38BRGlKKrE3FaUns/ndtbM4gRQLmaJj8oHj21Vtgyyy4iYW3xE18o18upf5nGOc7GwNQMS3E5+R
bU40uVqyuq98OP4+zLYIQsza9hEo4K6QASnog6fwYHZfW2oa0JfNY/1wj9OcP/nnKOAoHL/WNQxz
RJem34204JAFCwH8NIABvzD5FqUhZPOvmt9XrVlY4L2VrPdgIuUhI93ykWQtYgdfGgLTu57a8xYf
A1uDE0UoTVxkMBz9bPLaNVGS3V7oECK5T8oolIXRogzvOVZOo0/gr9yopVQWCBJajtPaQ7ig+TZZ
bKsjx1b2kOpkGzI9HvY1YO1z2ZEYIGcbYmJerl8fHm2s40t3DrR2zxmAJg5tPQT+/zp7GAN38VLe
I2sbsUzCFlFAQmz0BRyvinp3nOxdWXUv9EM/ndEOkRXPkGN//GzmhjUU9S1OBofgbJTUx2NJ33j+
OYcVlg9RighROojMydiND+bQezULLzWfyM2tzC3nvPrfm6WcDDZcL76rLRMvltR51NVKbaI92Bxr
zecXR0D7daTHoxDDG8VtZJj7Pow0uYQfo+M3dVa6AWsuK29Gbenzja4i8c6W3BmBkbDQFCLsjrF4
FYj0fYTT3WIzlSISYO2UKEgW844fxVu2mguPy8qFHCgx1bptcw+wQlCKLn/UtZ6DTxxqn5kE1hrI
eN1OlZWpMOQLGuf6oPw4tadfBbvylL9HO54PD6+IU1mKHUsvX0n4Mx2zEr+bxbzQhXnAveNBZH4c
bLVmK0bv1hoZwX7Qd/74e63A77fT150bUPSmuJbSBOZQa4bWqD/YMqMIIkUfxA3HEtX8/WGRWnBj
GW8+VgpnZZ7uBEaoEaY1wk3D/HQQRNLppqHAKvymXdf+TnHPkWOPHDJSDO/SwKYd0KW04WCD4Nym
aLvDGMe7cahgFUp/ySGtTf1IvZ7hGjdm5vWtFuOOtgTK5eFwrJLz7gwL2FbkczltbPqrt5aors4M
N+DKFrim+3hsLL7dgS8C8Mvt+HwzIw8fayx1GIg5VchWt+kJ9vVyRW19qhX9weI3Pm8Kb9uTj0o2
g0cKACl7bmVnA5qMdShxuknsIGka24Q19WjQbYMoo8SgxYSt4oOjj2R9JNWRyERTNSQAE7aSz8gj
FtiaG6+ui2OizLroMjxNeK5RDipBjyFVYw1pCnfwLIbAnqh6LoV00gLXPItoKFOom02OK/trsY1I
oaCBAV9I70TitoM/FluhMasy5Q+NhflhqtCbQ27w3CypWJf8ct7/6HOryS6zqOVk824f9tr8u4MU
gtB15eArPb+UMpU83VXw56+I8JMEPvp9qn9G6+lXFK7hCvy564aOMyxBi3PYc8hyXOvlGPUdu4NS
KppR/jhJ/LThvZOA8Gja1O43W+KSeqbTYzIvhKD44T1yHpT7sg1wjT+gYqPVYqjre+25eLl/mrvl
VeJxJcpm1hiDas7OT3FdaBMBSFzAzXtc6elQcLZPo821FtEe+DhlcKZaxd4Z1B8mDlUJbECwadT6
HjoC4WU15JNKCZwgq97GiLmzCvuBom567VnUbor6W5icfdW7NRoT+NIz+8WrFDDE71a7rT3etArY
i831noHh94wWvcuOts8yUB+c0QNr2MH/dhJfsiS6DuYc1DUlHwzH6GlAMf68TbbUErjzkVUCuR5Y
VGfA6lW6yzf20NZ8S8Gj+gu5IEshwc2C7vk+sYhRGyJ+gEBdkHU4ZdWPFGNV84lfVpE0BtigCwPS
PT3XZBFnCC5h94UxJOuRQmfA7EAZWjmd5Pozlr1YAXD+STYhL0PA8meH4/0ydjaBpItWpKjG3AmK
Zadh4MMjxrY9vZAMt9YiBiCTp61P6ltCcJoDn98BtKFVAqpYOD8nJFuOs5g7l5v8e3q/gCx59quX
rRryY2GpMcU30pqSC8Tz87AZSCQINSbUGy4yVVE0OPDOx0ICvRoU/OpbtyslYsBoEaQlYGuYD1ul
ZyArP+AXuOd3ELqg296q+9ycWdVoUv7fTnxuHp1ztSiX0wfxaWMIbtXJj5LNwYz6q8FZt2cyMlcN
y/IDQhWdWUcGIAok6i5JunXaItkkLIidFADqL2B7LP8mf4p8k9MgncE1pTKVOwUaEfEKPyuYXCsj
T4sd+Mr6cnMgVF95DBPT7TQUxTlA8GMurVEduaAzDGidBwT3XE7xqVnMW2wkecWLj7fFZAPOxohj
cUNOKyqj1TwprtxvbpeWW399yn0jAs2xLjCJz4/AFZ5ftXk6DrPtTZyo0GtVxLB7mcPiLG7mUnqO
zAn7vIJO6nNttq9bske+FckYZNJspHXQ4annhGmG9WoFnLnIZMV/Xwg07VAhYIsAl//+O5cy4t5J
U17KYNNM8bN8IjRXffj4rQR3O8s0eqLpatDWRAmFsler2zsJBcCsdAqtrDBvfCLWtWd6vviTBSzX
nUVcOoksgzWfoXVYDiXSJMBrXBFDE/3rcXCghKyqWG/h/MpVQ/8Y15iwX4KMYh7jyyc35czOX2FZ
EqVpAjEcHnIz/pZRpyLUjBOICfnFnlfhQnDKGWxaiTQ1X6D3C/ryGgN9vgFhPxMXzvEQLXEvZP4R
qzQDAgVv8n0Ydx4gNJYWLaWVVVY5Qty7eKoQN9sQL1Cp3UOgN5W0ojsJrYqPpfg8EGiVGm1HzG1V
syjOUj4rxc5K4RNWLQqa1JS71yOG2zssSuYTFzOxic8LQ8T0mBfMB5pVZExslJ3vbJbokC97o0N1
m9WOSrMnvPi4W002K0iOwezthn8I0FFhcU89EXngpuMY8Rd6JGFhrZ2yE42sk2NUwnBhQgabPJo7
uPGkqytobxW0pFo0TKGfCXiOYuHV6nTfTvoktMa4Zh1+keURlpgb0kXomum+BVVF1HlEUl+xcCbM
SMHHflrFq/oWdGlkA4S3MF/HtTK+IO8zJZEp02LoeDYNrd59PJIo3fBN+i/i3S9W4N1SJjkjPQkD
Cr/HbKG54GjV26vBLPTsEJF942RqQaW2Rgot9IUHD+O8OG7q4NAjqsxV7TKB3OWNg4RRevKOyvaA
PDB4HzHXBp4tKK1O6s2WEmrVJU9AU7dwOVdSOjMBGnr6SfV1gSAWMB9l5vv1s9V0qJeUt7gn5VM7
fYNSHJCqeLi84DAUj/n1JTlOrWBl56pQo+qcLr3CogE0PVfUBuPawBQABkOFi/dXy53p09ygsOy7
OSXmgZ1Rv7RouwmVtXAUX9gV+UKoBUBagsMtzADGYXA7mYUkVfE1DFR6r3qhfQYxuu0qWeP48qTd
6mKGW2necpDttihgSgdjLCBxYG2trm5XfxwTJ4HhY4PjvLAEbGHlMYmx656AJqZ8o1fQ/9tDZGrJ
jOfHpblPTmTwUDTYXnSkLFmc/VZHS+RPmsOWvrT4NMms17nKOxiLOet5zYbU+4QiSWIhV+TJJv0S
FS3fYa5FAX6bjXO5EDZ7IiborAoYLpo234EAc1iMFrciAtcG21EWMJiR2xbTD7Sd0Js8fIeOddcP
WSgm8aqge+WsUjNV5QV5D4kJc3vD9O/l0gP4ZKVTdoH9wzjBARRxo6np4V1/+NjF0oHGB9VQ8ezu
9AwJvPkJefCrTWLDM5kXP6vqQM5K52NvDjYe3XZKB/miwgNGU+yZBzqRMd81pBAkqN126gnUEqaA
fSec2Hz2EcLYyZxOtnCkB8SqJnoe3bt/A9UWgGDL3VJzH/H0vg1wSy80YMoZ04VW7T9Axp5nWTHZ
beRy+QaoV15PA2ONc3emnUYc9O3GR1tUZGf1lJtNRGz//Is4mSpCLCQeM/eKOH0vQ+w5t8MF7QkX
S9LxQu3m7DhVfQElCAdwU8G5pBblHkg8Ybt2Ci3lFc6281d3lzcPlwKeMG4u8MYGnMrrNV/oC5bx
pLoM06GTv8P3Umf6cKLuli6bH9FrFeSUD6GXpyAFDnE2WAJciLDV4hSEISC3Cyh3rDeHORij5VUk
wy7YkP1XE/R7vJ5c2jouVatv0aahfKIKhQPenwpG83oKeQGwZWz89X1HnR/woWHRASNBzREAV+Xb
y1LGAgEyEdNXTyaVVGqklres8wZIJcXwMMihktHglNFp1qgwbyD6SpyrEVavdiu8VnaFOLwHOSa+
DxC+deldybG2qb6UEYqjEFeyn8nXXt7LGDllN2k1r96krujxkJfLyZH3V64kDWA+L7H3dZOYaXz2
D3Fme1tWwO7WqjHmaiXQsEl4q8tng69fTzLwg62Q51A3/sXqO2uXsCngSz8unM6CQJyTqCxfYo9m
DDsTP95kmCyJCx5Tos8diORbXPPc9KMNh4auVH3wUYCREjGaj5QXqDWwGYH6sHx240mIpqDiarJC
5rYnBNvgxJyiiJVKKS5jUzOq4xRgyqLnXROm8gWhaOqQqv+lRAPKQglNEvb4y57QD6ai5VuKYTmu
P2If9f4SIprRpEuTDJUhECLPaSb+WpCXNE9tmM9Ml1hUMyBuZZHBm5BNxzoabnT6B/0/EC6j2y+l
EjV9qFkpCoPvZHRl+9BZPtHnQAEZIsNctgrMGRrNsFLiyvCisRE7BaTg3vOUpXNL+fjvr/vHm3gq
eZR4It0VGRxevWq6NNWHMjINNE7Ex3vgA97NahtL9/r6wHWVZjU1V3sz8QyBT7J8K5coyE1jRTZs
gqc3G6qjS/nlbfgEQTMb9UcjyUCIayV9K25B+Y+HkPfZamqAQCrtW2PuzgjV1vwPqY2HPpK6dQKW
V2T20UOfgMYTwP1+sA4IpRQwDSYcsVInjYQ5PA0DTxSPbqKRkENX5/L/9i8BS7xt4kKQUCyCtIln
d3SAb/mMJ0JZj/vkJDYnLH9hiXLmToYn+Ezcv4Y9bKeZPkv2UVmKys4REoDD5wyA8Z8GfjLXpFpA
LV2ruG9XFNrWudKng+uBsVBdxWx22+XYSAow+W2tW1WubAg5WX8oGMbzmAnMhlJ0ibFYuAgu8z+D
o4eh+MY7HZ2n3DbSLLulMxtYuMrsaolN7CZiB3yAVKCDeM4uiaUB9AI9uZuaBghUxeKbHdh7ISrr
2tpjxyNt+qVB4hSCMO7Wl4d8OLfl0jCZqZlQHD6j216mCU8bFgH8Q+EsAX2Nx78numCVpUqPHTE9
aG19Nq2/2PlFL+yj10cM0ehCdeJgp+UUgoiuAxo1mdOAbJPuSor5ZWgMDtUup74dqIbtJK309FeA
/Zkcp0i/ZfubUTvRXdVKPboEPoZz318x9NNLjSpoM4Dl3Bql9EQRTEKH1Y0PIpgJUJwOk7SIA3YT
jlaIso/nJFBXgYy4QUmBGn5CrbdjCaCnA2GccL/f3nR9e5DID5/jYx9wZ+qL5ltEactWlADAnC5u
YB30UqOvSK5+TXrzHgZclXNPt97hZ7nP2NmrpXqi2hgvhn7rWBzxb2xG8aqlLAB8O3XBQemk08mP
QcOqh6DdWXwCfnvJdHh9ZjVgR8gfNZrzo6bXcF3KQWTUboDgs2QfImYt2ObauNxeAIeXV9rX2TlR
xCH5jaB/zpi1ian7Pxf0Nh88j7MLF69dOZJtAiwcAnm4NZhhKM63naPTORP939hA7WW1euF9SxX6
8skwHaaFoMo9yuY1sHAearl/liA8iEOhJAP2C8GPRHOvcu0ffQvRzxim9rSmuIANMraj1sXknLhb
7Gil2VyphsMtVLLCyrQUH3WaA1rm0ge/aotPQNR4avfQtzsq/BMwE8y0D0b7veTl+Zd02+Zq/MfK
yxk/uvqBfKbr4kyk6SmgrO3suCzhhxecd7C/L4+vuEl6w3CogskzN+FdYYd2SnkYpR3HngSxCxYb
5RX7zHD8gwfHNssSRy6u/u77or3ia1FrHzbhQXaqZsPAaOgEY5/D28LuAuon+4VBnRO15cGtxY6Z
dqG9HfLX/KgbP1DNJpZ4YP6HvviZx4PygEfCzMfqaxwt0K8QWgXYBPWtJ9hZ9U0JrpRYo/CVGEws
JTdxRlhRJc7+cU3oosMXrsQDgFtnfC+9JBkSbxE+RSTxUGjReFm+rEeRU3zeD3MiLz0sHCXuozuX
s8PmP/GFD83IRIFCOIe7hFrWrAX7zd/FWo46hDfWRjzUrYHf9AyszHqpD9YQ9HlDb6SrTN8w3vWp
4Py1K0pc898OerSzFF+mMXl0HRLXXTl7pLII9nvApoDC/TM3ueLTGvJz9NUPitW+bdKSMq/wPAax
A3n39D6nyrNzCqqTUWYQNAswSNJ0GoaMn93JCJSHc0D6ya1Hjl68ylgPlAM6iq8oSq69Z0aTLamT
sCHJ1XP3Ag4ug5puoJcoWH2CTQUgVkosLWo7mzsZsjA4CurL0fvwmF+Nwb1aXSOOY+QV3wMEIlD/
uowObnOxGOrqPap/Yyc2eC3aFVTvq7GcnH3QNcaanoAJZ6Y+tHGi3QPuGbWewebac5STaEzOHQ9j
ddKWgE6XaKyxygiI3t2fvrhxf9aBQri2ps5FzwYzk9M4IESAYy7kDVN+QNdDHYki0BgoK96LD23g
8x4nPasHWS0YWHooDw2JSCGSGPL8zVT7Pu1T3/Vfavwu9gxmZOIbHtHVz9PAX6uGHH4+Qt4MRtI9
3zE9hICntIJg8QjqJcjqNoTuknUUgz1D+CRIiCznvwZX1Dw7UMhEfvLDyZWO8nW4NRvbp2Zw7kgx
QE7viCGoy2zr++nlNUIB/6mbKAi0QNWUbe4WVdWdXqon+Vcm4O9UhJgUIxExRWM5ySNJZZ5fFtkA
9xz5pV4Eegk/oPnGseqo6hAFsMNibdjvGbkZtj4mrFNOeN4fKcsiMVe6Sp0e0QdiUtVARRH08ChB
8sYDiI0n/WY9Ex8O3/1QbONhP/G6Wb+VF/GZtRr+SYqcQhyDlyOtZ4YCPpxP0Pt9015ZU6hes78j
X/CNts+WRdk02t5GezRV0JN1/aQI+Vdgr6drK1UmH5VrVAmWhv3Y5OM05D88h/oz4BNGdc5HCHhF
g2ozwgvpcBWxAwq2mTxSGDwVOCBRNWuYWffRoowtz7cNFohzjjrLAoUoWfQAgO+SVu9+ihRTbWQG
h6nVzvxkRONds8KwWRlR8FPg3mTUMcyXRlg1fmIVNzinaZsn1AdHciWbnnHdbKTpIBjqYxlqwuuH
SX/UVcbyMrpWMVywfMFe1AOcF6S5b41DtiPtkYCsKx5sSbocZsZAXugcZPn39KLevruPYdAvCBzr
aJZKbIWHicsbUZ4F+/31kcANfRc5tcsmk5DfuAg87/PktIxzfkLYrNCIdFHU9nJ9Tvt4eWheZiSi
mcCmgdpKQp/+IUDSVrbyIAT9aXQCAqs0rIv6+3f3+fCmgXAniFZlOmBdvvqH5p0udQ8I0bq3NDpY
30pKBWXOHysCoJre2G4uMAef9EX4jwPnQxh98thevT8HEubH4MiRdkXxazcRcyuQZ7O/hg+toREm
g/4bVmvH9/1Lf6PUvAJHeCT5rZyt5i+O0AVgx+LoDH2wtCh8pUQDi/ISW9Ar1UOm5V9qMfAwKnI2
WWLGsvgAXh+uFl0y15te5lMTsi8nc8+MSe5+ONoaKh2wdZZ6k8YBkLL1Ow64By0sWNcBK4CoJwIN
F8V65wL86WrPip/4j3O8FMBgLjVLQIlaGu84LQJWPa/NQ2hax4+OhayFYKFIezsGA+rYqmWjR6kF
BfgrjFWaGRLkVmCvw+LpxqFA4ETQIDf+aXwVYNtZgai2q/kQ84bXqzsSNGe3Gccr+v153lD5J6BN
pZU75Ewxn9Wo1DGV70v2PwRHNu5il3tCBXL05oX8syvxOeUL04QtxiF37t8P8gaRJveuFzBoaeK/
XXKfuxANt8x0WMs51nw8MY0zZb3lIodi0JQJ9rcpWFC8/atqId+sVKmUsfwUp439c6OfNSDKrp1w
ufaPgf6sV+x1KiQa4z1jA6BeUyAXDEmU2qgbCj+xZ5WkUvU8lWMh1RBKnAea245tVgVcK90BS/x6
dIL+O+ktRRCqz7nArG+n+YPZXwqZFFdWgG4nvyNbW4qNbHI1W+5EjmOv1SyGGd5oFp21DnLSFSI+
kG6pILRaM/tWVqBni10xMXAV7OHmS5AW/1WQzsjlcmR5JDh+Tj4aZRQXXSyY0h/KqsfDhvGNYxl0
nRUZq2hsXpjesOoEMENKvydlSwerYxHeRrGxShvxQBvEkKBy5Ia0YdKKRC/GeRFWLgmGUgGWzJfd
l6UhMao0kZqJKmGaix9d7koWZ6BHiuWoGGAs5Bgj0oRtRD0v3jS3gmSkYQWrmd+68fV2dQJ4Lnyg
NpajA3h8RF/tgTbfN6KYyqNj8Kl1Sfp+K3aQWwnRuts1K4wxV/rnHxZmiUIBa+wmVfKq/dMFbbir
/u8Cu9mkPDiXr5pQjO3T8zas+ZqJmyOUN7ojZM2CC/COZi9GhxsG39g+61kuLUPv4kKAIAhO2OhF
c+nZQABHPmPvqsZQiuCGcdn6z/t7fmiKCM90YdNNuDSFpm5PV4erMydjoSpMscHX6v8CMWyKMQF+
PnVACT8hgGOxLvITN/iVNHMvTJ4VNKa79yilWBEI8BPnYuY/1kFZYv/YYln77hTqT8naqeGYmQKf
Up1WLvgXGw2ZzY5qsFQpOnfafVWxpurjkRySZzUdhq0V7BbJSExXnMn7rZMHYLM2JRJokINfXEi1
5XEjbtCQxDpqsFgpRrJv0FJhHn6UxW7m8e1ffFnctbHWJ6mqEbQ/LMv1auaBZGhu7AD1YsvQp+Ps
uSUMmqNvyWDs9V5ikgi1qFUXG7IiMlmzt6wRHMVUSHMzGaoizZRlaCZrUxEBLVPCEf28xRlluJFK
Au7E0ye6GFL5q29gUL/NIALBrIaQdZMJx2SStg/avBrC0+ltS3pABx1JrK8Z2Fjq8Ns8ZeTyYAHL
fPoAA876on11CuydqkcERkBVZq38B7+/HdHBi7FY9tCd6AwMkfH2OTH8CdykTxKDSUbn4bEuNZkT
h4dYv8E+a7+wex4wmWZ+w9uIMZkCTauSyGIVdjG+qjBpk7K0I4krVE3Yjlvg6+7jXaBt1kwxW4/P
3htgy/n1vRd1m321V4CNXINru/RLcXEVdRbHC3aiPPPepIcFfT1k735Ig6NmzHNAx2ZK3WSQ5gRI
z3tiAuixVx7tKNINDicgj7X8ptwvoRroEHf4hUbNDb0hEJMFyu/m150Kd8A4ePtSsQbahapM33zv
wE97jGhrxV9EoOp84oR1kU+eyAAO7/1zqeDp91xIxFugKSaqf/8icyi+NoECuEcVMxoTfeMzp2eW
0S4iDDqsBOTUwTMIiY0CNC6wVxq9B5q587Hx8uaOoIZ0pTt9D9EhaOQmcbKhkOcLNkFP1LwJHI00
S9fPbDQAcgRmc7T2WhPq/nP5MtTHeZ0MkYN+BJEUpIM5CnQUx3RuLlFp0bIsBCPw2z+57GSovOK8
B/EVwn9tNuMOLpdN8oxAQJmn6BhKDFlvN5FoMcG8BDAYj6Ji8hH964eshWnAHzxBJ/pKrwP0at4j
tmUETI61HKUhHzQq4tw6RvMS947yOBRIbPfO8HQH8yC0x7jw24PsMPieQmapNHLq5labJA/E7Beb
vfZs2Cv3e6EQa9e2l/W/9xxYJmsRjVOnhxtP9RKxbDE2rZWdjPMouX2+I42ZguF2YGl3aSg5xsgt
titY1ryFVUi1CcXFh/yCIffveAHurp42pBnDc82e5xcDgzkY7PAK7Hw/ifuqi2nU6FeZghSyvYSX
JKDF5gOfU0Curn3xKo1NaLEqKSQRe1miacDjNHFRFrwAt/M1M7RaWQf0dBTHTk2y7JwqRoP4JKTr
usKZDoRxzLRflBeeKbNS4JjX4WOPzzqXRw+00jSvRLYp4dsNRnxElUlLb+93kMAz3SD1k8WWsl+f
6SEzhclaMsZXr7ZS8M2ZfNkAX+tqeJ9N1P9pV5oYfwamnGzifjxTLNmdA0adgBnsQWHkjg/Jta5t
8XsUh9UhPCKkhLZyZg/o3Atl0QTohVyAVaeBlW8MNinPdDkwMP9pV9rGzpHeoJGt7/VCZoTne/2b
INc3tINZVYT+eMezXqXpo8qZB/Gk814Za/jLxeTj4WF790cJvn1qMgFa7AGLXrwFfx6DqzNxS8+q
5cEyoXmX3LdHUAHmO6N1MpwVGi9qzxlyb5Vkh5tKzo7ErH2Bk4y4lukBcvuJNLML+K97QNhPtcTQ
9ILrMFkxVa0o9Mm1FIqOTkeOy/1JSc9g8Gwj8r2WqlVth5J52CvNBOQC4zNzUBTh3fkqFTgOtfFt
EdiJ0wzFxn603pSVNyd3Jhj6nl2QNkIluxwoUJRMRLPEMdzBspyTPXSX4m/0FocUwT8mGeVFb16d
cb2TwKsuq3fXLluHIRb32oIRYoBpnXY7U/iaDNeGICY1njFFrRMk4iYFDzkj4maf1e4j+lyX0q3i
3v5GosDfAkv6eq0viHmdh8gQT0E9UN0NAmfqTpYlA5/l31XFyITty+40jb+Q/rxtmJzrt3VBRYI7
yGkFdSSXwMxlr7d02L8njIiw+nR0HjExNOhjP4iZTxG/SKM8wOaoBlLR1Roeon67AOQVVagg4MaM
2uo5tnQ+9fZWpczD/7SSsPDrdFo6ejaqNENtX/zQLJVVRcORfc5sjdFOfYmpstiZnZbC7hcafOrr
2bLTJcmmxHfQeEdmbFo5fSzcTGH+fKwaVVAwny/bwXNb0v94iCVvAxYH1JCMdoqu1WhZmliwQgvP
t9Eqh7+dHlQUCrfMWH54KztSf0jLnHrYK3csePprDIEUBIKecVUNQNVS8SGGqm/E4ftpvBlFHVzA
pUlNCJt+0S51ZuS8Dc/ySE11BEnkW2DIXFUWxRYDSaIvAeNi4rqclpzT103kFLalsq/JKVULNgwg
ZXATCxoRV1ycmQL/QNLwpTeGQw8s5LTxLFbN+yA2uFwYNShsII/zEzUIxZ4dryO6UBIWJrhYQgG/
zUu+m5t5Xxyvqrq7zPlOvtShac1Nulimab9D1DbX8IgExNjBec9vSqrV7ttO6EuqAjnLI8H752BC
wYcJg26W+vjaCg6Up5cN0xRACwy/NoPf9Jh7/YtO2+DHRG47Y4FU7oYNydXZZDs6Cgfy5VI+odhK
QJiqt1EXFbBkQaM4Yg/qwax/a9vTEzvdz5jfLCXCUDZyv5Ha1MZcUwcCJWcqWFw7guxcESkjsf6h
vHkFu6uTdKzyX7LZEMBzq4pFsSUpPk5fgIPsewsGQU64Eoj6Hm20WLIQ2V/Xcp6jCcgSkXXqrex1
tkj9rnMv2cy4WcyX3/ce160L3pua05XyFgs2u8W5q2NKo0iqcsAOPs+T18jTVMPGHPIAFejKyP/K
ndtz7tPdnVvhfG9nzn8dxb+y5IYHSNJ8mJDCIh+4sZ5k8aORkIBc6LiAafvHR7s5LkXo6NuPgjA0
re2ExlmfspaDQpaVElF0RlyEASGoLHHRdEki723m0lKTuvNpfMG3NsGh85ePhC1+kcSmgESvjUrB
OJfeCii3syKn1Zhh3phAubrNL/x34yRhKKZctigQLwsu3Csy9VlkCLavfLWNL0O7c/47Zl7qTVdZ
+9lnubXmWGfVAmul0Q3OxeUyszmEHHXcXWISRmJVAf5qW8tY68ewcJdPQi6BcsQEsjzItgWCgu1Y
2/GyMogyBaB+eEk5NOMskaGtdehshAkh/HcQXVXRFoBvrHTmuKN1Y0h7CUfJNMVISrGTmom70BEG
XnSqyARTR5fb9jd/PPrYwUDjRqAlVip59e1UaDQ6UL9TQycfPL3esoD4dKTGvSaL9Jm36336s83g
lNjmC8QYAJnpiOLN0MQdCoqw1PavTGVHaypSNbP66136umLzUmYRdTpdX9kMHEWH6BjWkMCbT4HK
Z2FGVlBQn6sB9NtcrSOo6qFgVbdSo6pH7OeRF6u/mtwfiO6WNN8OvW7oSaBrkzdY44AgpOQUAOdF
rhgMIlWUZH6Cne6qfaCN0qKYDUHiOZiss4uCVWRmFxSPj5Hlw/fatOU4erA3h30OtreybVnuHZQs
j4kXLVaJM0Y96nhYygOh08xNa+bo1Ho1wA9Fq7HrDtYQK4pvHgYuh/d8cL+JjFW2ms3WQEXm0Ulc
N5HFG5x7yBrrsbL2qHMTWBYrPA1sVpMghetK6E+7ulh7N342jOyFtMEIGFx9YluyVG/D/nbSXbXY
nLgWilOIRhPXigKfxvNvLj/qwONNVNHMuz35DRjWs7+P1RzHkjFwcyrIUrhB68Lk3QgOBJSIPjKj
0BVwayZVBrzkCqKTlwYAgLtWyQivGLsF7mr/SqeVWaFu1bibsDKV8K8SlbICHbGVQ/tmhzmjOD7k
c/iqGZzEchwR6I5tpE4vaHUmrpGzey3e/3w251ABUwfqBQQKMzVpOTvRGWCq6HCJdNWwniEg3Vr6
QOzrqlf54X91Y1pZaqOzxbKXg/EnYy0iHQBeVNAiMuBhump1FsIBMjaacbGk9TV7OamKL3hcXV/l
Ntl/b/jjw01P1Yo/4SbDFttKVuZogpt525nskH+AqvNuOSlzwqUXVZrvW4gPgc7exa6OkIl5vBqF
dhVnUEXRJ3P4YaEUku4MwNHXPE2DN2AhGYvgplxX2x6knoY8mn3K3MhqSsCUSobav2FzaWTA5ZJf
nCQZDZ3bfF43Rxc7AJ3l0dy1+6MXK/1v7xouf9t24m68GPKyFWQlaoF/Di3kYvSvY2Ju4U1evsSr
n+Ff4Pvp2ESPt1edrbtuAt60H+SeBAy5CrA7X/m3ejlV9fREwARTeW460+Fhv9C57Qf0ncNPuzgh
6KPsEbvIpql2SNl5/oXusEDtsxlKQg5ApgdZadXYAOv8vr110FP51QB72oUg+mHBqZzDU7IoxHLx
kPM4FA/8VfYELKrsCQCX/Ru49vw2gIGKELrU4ZDvMMFomQdVsOZ1j4RKP+xfYc3JeYcnntcjwk4f
qdud3vxRRrLCH+m1nVcWhIN7whW9xSg7qUDqseYO7Rr5s8mzY5p0ZrytaV7yKeYTvUy9WnhIBXHV
bB5vE5h+YtFmxgvdNXS6yddFlTVvJtusuX2XSESyTlbyzvHvvv6jm1RkwViRF8eAe1CW/qqIbYf6
Pfy1njus/vUb9hH3fMwRAtsB980jWK8mkJNV4oRDGv3hCqtqfD6RO+ynnVVGQZWv5vmhJqEj1tYe
rLYDyLAix/+7jY2QlpLcNP4gQCxMloc/q/WEt8ooCG8OQjawPpdgeIWDdig8JuucOi369Ac/6Sio
l4k2W6bUUQ/yioRbvNQMPtZKu5Zu4RqbJ/KFDDwzD3X+AGJoxOpyiovzZB9z8v8nln4je8mnVrYx
+kTkOBH67SSV6ngQDCJLSAjy6+ITUZHc7Z0q9HWomiGXxmtvvLc/6Wgrlj93VO9xl1LSe9PNLNgB
qHDVppT69T8O7qVzdu7A1pLyE5iBPgAmMJ0dg98YV/gVJZd4LvhtDQpydzXrt3q01Gi60lFCvjTk
AR+/WjqrpAiKrJEFwwjEew2sRsr7n5c/2/X7wDvxw7hagMeZp3OTQsN7r1qb/zFqXEl5jDutouU5
cTUT8ZFU+aSN3YLxqQGU1pi3up6LFY6bqC5aPQpyydni+LP3icmperZW/YfXHzaArMpKJxcWC5pq
VmbiMtLdu5NPI6XB7HYoYVKqHvHeSJrQTOSJxusYfW1Ue8aWQgD6Wu4xkVN3SsybjLZsFCO6mz5T
Gm8qRihNk0GIxHLRVS6cubLmQO6LSuEynVfwJoCmryksMiHFYQOLLiZ8U8rN8Xt9ALeFfhi9LDVV
5ffS4qXYEXt89v0d14CM31fuhqBLNfva5KhFfQD+lF1UO85UzzSWNoPQnUP1hV34AZH6f9Zqpzgj
/x8F1sPMK0GNvgvYy0XylNlNnQa/WnAN+9vzRk4HB/J78+fUQhpk0s/DVeittPdlIaLDjFWnualY
o0PFt6tW8uhV6HehxWV2caia05L+RucM6Oct/UbElQ8h/M7+NtV1J0JMn7M3UYKcCmle5a42TI7X
Qq8gJcStTMy5PxGEplcrF/pOMm0gWwEOW7EolkI8AgjpVgInoKhaySAa2Ke9oRM92TPvfGr5DLP2
PC1KKm5NTfybeOzyxhCKlgezF82/fU2bJQ9LQbBvu8H1twmFERB9OGquDSBKxeTPYQ8pJDNF1OXo
GznCKewzsXh2GeOvDR/eiX+xuUb5rEiHckP+6IBFipRpAKzxBoCtL0scwBvocCzNfkbCGxXJqQmX
eOzjVCOX6COaQRGAW3xVQKWODFI1Jn/zrIlZhGZlw35Np0lkELzyQT3bHoIS8HfI9FsuPKGGLnl4
SvMsnmsVdSyoYuVdWtqPhw6cTSUGmhH6/o9MiK2tidvhum7Q0sWMdIMaP/nl4791teyC7VY/ozZH
U7eD1sfDi4pLIpWMRHNTlyW0V6pme9/P9pDLRke3tT1JN8hne28sMwSGNEDUpQAfnnHTdDJR0iAy
/0VEY+gEY4Gsy87u4d98HnoGIKeRsM94wnxgKlkvIxA24ss5+TtxZtnBvTWGTTIsvF0gRq5qc7mz
OltDcQm6xHZUvvIXUe2X4z20udufuj1cfyuPgPCkVOcAIYAaHeBPyeDZcEL1Z6VG9WAGs3zxtgo5
P6rk/HsElZkfFUcpKTnVXYB5knCb/XplaDxcoPnBnHLc49xRxd/NwIeMMIbOPWbWN2oMlFiVX9/5
ElV5OuSW2H+ZlmNBqLivOnSrGfOBzSBqlQ2ROymNBt+itJ+2xgB8cVq+UwIwkuYJOOngYOycTAM2
xj7uTAnAWh/HoIDU9/smgn40UHSIqWXKlpEIM2bDXnqlpwJylbUQ84xozNi3DfJUO3RuCftD/V8L
SsENf4ueRkCwebmr0iyWkdnehLqoRU2PR+vL5La3V2RUrV0i3a2MCotmQ3Pb6KyfTx7FNXLMNBWR
H4W1Wezh9cgrMOE9GVH6YlON+3rdrnxPHMdh3voFbJQVMBtRb8oD+iQkmnNrd/M/yqFUfxlUn/XJ
IC5muf0Y/TPCz40RpDCDlfqkLU4ojYbBMUcwDxMzHZ7VBHqq9cDwT+HyL7fJ0HB7XMQD4YGJuHF3
U9JiUlgnB+ijxoy3vymkNBPaJjqg258w1C6ZypibkahEIMkoX8uMkByz+gMMTTy2O6fR0ym8hCcW
dc6oIvGE+a+OTZPv4NOVXhBdZq86pvyPq8Dp2yvT7WpIZ5j0ykx1nQ/AkqCwMLTgMC86pqdrogDS
00mKGmK62M5Ah0YoC6Meby+8TvQSgMF3Zw+NCsuYqTs/QgHobn3vCSn4ECL7ATv/IhdTYLH9wQoo
A/7gLNLBfNhqTZQMA1mHAXu3+Bl0RpXjfNEKh1yIq02Wc8Q8VO9p0I2HoXnu5mAycIB7NsVAtt1J
ma6uBoqzWZ1ObL08s5iIupgZI+FqT+uhjrKS3bNnDKQFOPTzLFzgRcknUh4cfIuWdH7UtEu+xjXu
O3KAuo6igSPn6gWQCCGGPKK4sK/2UICMVVTKuRVcujktao21ZFMR5cge7Ha8RJGTd/nKPo5yitAu
2ZUUt5IqwfHdf6QsaAZapH6+8YfDQcwrAigg5HTh8gpWjmBm6cHg4Q9AwEAQzmFJHZ7BX9FRiFHS
437iJ9Bz4c3NeoaShPs3/WYCt03C04Nnq8p2aC9BsY8EGGBX+DZKEq1DbKvUNuRYYjHVCAUVydOz
z5gz68tUR6x3G5r4/CbOFrV/0jf3iDK44bVOHuuhtnsGTxjIdz8p9ZCF8/o6SXyXznqJDyd/FF6Z
Ox7I2yvdeqNA4KRSGOnu/BinYOzfS0wuXWhb+YC6fB2nvhlEcX5Tdk6Ap3hr98FzY8pDgtq+9CEr
Gh2HU6wdOa+DDL9falpK3Ad5nPSwqmJzjP1XIVryd2QwoRGsShXeLqOpIwm1IJtEqioiWDkhcJO7
bFlj66QNSFdbhSoc70ke9qBAm9AhHg7vzoTmJMOUHonFqrbyDIbykUi5pN77OXKtcSUm9mBqOy/e
coNr5ogsYDVncjhVBprRYmfCkNENJfB4skOAZsmQSWw7e1MrFVV9NdwHiawwmrBa62ADOfJJ4BNO
8+xNVmsVJ4BefVzePzHpaPHUQhFuGZAOPfaIDcJLfiwRVDMqZJA/95p3H1M9LXja4L/uKbgVrgIP
8AYtUXflMONTx2DCCJrcZlaOCWJCpsqNFm2T4PegAZapPr6hamMW3cmsmJvujickTUxjTOlmkzNE
EJTmgdVeINJ6pblJtAkjlHpvDSCd12PSnh2g7GIv1PgzKC1v4XnOZrRZX8bI92dVh4umLvMT+2bp
fMBGodhi79I9jKmvDbDZDjnyd2+X2r/eGg3SQYWfK2KKDiJbAcaNNwpbPbGmamKW43XopECYUXyt
biBfsZr4f6B+xSVFRvkh3jFWfqGblIK3G16NWDyYGdqQMrFf856jhm8vSq3UujG01cPBkzqU+8BT
UrWekMtyuV4NGarzNavsHMAsip9KB1cQvzsm3YRSpzxMpSAFNz2Sdm7tRVYFfseYj688tBoWsQp1
MjFtEPO/QNgU9KQM/mqnzWZFW0r3lYrVV3XhFhkLGZcfbwrLbNU1lc5NVzHLT+1xxqzYhy5yos3p
mSLpEQj1Mamss1k67DdGSEGjn2Yici+GG+KY6gANRs2fNHMaL6xVbbk3/Xlb2UBdjea5uogfXjk0
2j/Tfn7F39I5BZNvEiAJEK39bDWUA7VKPTLGqzpa0UZKIkLYOMzGHEAPufSBZ8uYFfx6z9TgGRAu
gZYJbQ/GQ0NUNg6Hhrhkfucr2e/0Wew9W93wtF+tJXIHs42zWH6cZ0K+kEq2fA8NLoLCD7TSl18c
rAxFuRUqQ6y5jFsPlb5x3t1tkkyLQvbcQ19bQPZkuST6jZ32mtztnZA74k0l+cAOa30LyQLoeLWX
umcF5JmEnNg4rGbn7KkDJIg7IJm5CvbbgPo22hhan3aRjxiKInblLTyW76og/XD2dqoIguJdl0XH
oh2Pztl9rYbbgLwfdr80MqhElgIurHkL+EjevSXI3T80tBuRTCVzq8FeqeTAd6dYDQ9YOhKUPIHA
KbM2SIgpF2iDSocFbDgkxrI1k39y4sabH3eNQ3sKzJm4s3vJq7Tvd3x8R3HQVBR1v0oWgFaXK8q7
PtK2wSTR3jmg3/jDeYKfXpVvnCbG8+zHM2pGZdakOQRdbfScw3DMfhEVeOglWUkiGkKYpWtzNrp2
wL3mVdu1cq6ZzFM8wW/NtAGCbK01UOhPbo07iKJlUOM/I1cO/3B7jlDdhkK15sYIcDLIe1rnvx0u
GQWjOqmLzLUQYUwzo1TvMRtGvWibFvLi+FfFbjCrJFV5W+KHjEVxNCgo3yCwXLoXWo4Wwd+IFcCw
kBN5aGc2iTd1W1ORtY8BDWQJ2StrxuQjZFrL74CDfOVirV4eaKcYRMcwJHW9uDikuH9eSKojPe6g
RhVAz9JevKwDmBxB9XaVhs8udOwWUXsYwAmV8SAR1btNHJvjRYCMb21OhG3AYVp8S7fuTw4ChcW0
LD7vi4jHZ2WFKiFmuMFBHysmAGJa50dtpypOFe2YSVtmPI0dLATfWyonPt/ndJUTUJVWaL2Cqodq
4mBiKFVkBnCEJaVvR6R6WCt8cOeKOn9idcIqci1RSw/T9kcCYTFqdCfhD3kPAa2OgSqmVTfhscsW
eEzu3O2qr/9KyPl2sRDs4SMq2H4Dw9cmxRREbV+D1oSnb0aloJIKWjSXAwC3O56Czphe5cP14vlJ
rtKY6hoSYYUBsOxYvjmzP95hf3j9EaYt0pY68ZK5BonggmYES5aRh7FTRmCnZGAgoDqqojFVd2BM
xdUP6rgwp8Pr/D2cRsay9M3CKErRu6MNTxvi+ZeDyNdOqRXl6OXraaRbIQjK6CU/PZIcpH2JDXR4
Kj1bTSp5iLDbzESaRkgBTai6Ss2knqsOdRWfDQappgKF8zGDqvWUoq+hKSIHTBKmNPg+llDK8a3N
P5duOxR9//Y8mwn/9ouMWq0L+HNGITvy0R4Lb9V/hYpyqTDp0buvWBYiLdEWoHGYUwEnboiXbecZ
2KRTZVYdiOemsAdfubqpOqhyPmYiZXnujhFMRwLY5NiGavtihdPbs46qGXk+p0WOxuxfy9HBH9id
BIolBNPaK8fwdap8NkGWGkcT++r4jM5BLgpSJa20NSkA1hiyH96wl5X9oQ78C9U25XgZ3dbeObCH
z/VR3ZklCFWn2yFasjIG2PZoWYmhCHKvCzF5jrDNMhXmub/vLlUEsOd1Nctm/oOXU4VIWT/uF92j
gi+SBwNTZpXAIm3NT1ZkJR4TQO3oW/0BbR8qqufFOVaw7FSHdKeRwy8Rk8SUP2rraKCKv59jGCpD
WIoweydEXEbYj1jKE4NRTZYuZJoUIec+koVU0Z81SV4L+qJqf53B2WtvGyNPcl9lyKFuQB18Ht31
nREgrFoIw9l3TcG2686xI6c9prsskoFR9mDtK3usu2KB6pHb1VeyWdCcr4lD7/QxysLQkEURsmWS
QOy3cm4i6x3gagQxseixGhM/85VgcDY0segasRi7k33NxIiSErYVJQPrwvqVO6l2f2Ft6Ue8SgsB
nOCcOt2gwce77CCyP0pDm5pC00APIxzunhZLJmhUStal6uwAHMplfpWBjvBtglnIA44YFQCJPRpl
4zPFNOpWPxEts4+ztyahEdNjtl1RBeP6A3DTVXMHX1iRLjOgdQcd97eFC+3foFqnEiZ+HmFnim8A
qmp6TNell+3R24zdWuUBYIBO/LFsCqHm94o8SPVZVkpopS7mkIWoqDJmGryaMhloqEsLBevQ4tXZ
VZStjcn+rP7VKJ5fG/15oTSlKyNpq0av3IiqQL224ebKdPM0OcHHZbzVkhLHkfnKzBxsf8KTK70q
nvys/SRn5cJpZ1re0TKCrydluiJVjjZ1YlrTjRhoZolqvBoxF4XU5UQTbYY73Q8LTN/zm12b+JKx
tpDX1nKFbwqeQoETFsWhav644kZ5YEUWNNX+QVEliMcZKwsEXRz+lZeUH9gBkY2JEr2g2rVTLEZs
sfFqt4ff6KaWAUnA+h7wr6YdjfYFtfrnfB/sHCMuja5CFxXtnsZKqtzoF0vX+1SxGsy1Tj0WFOff
CP1J+h/++Qwpn24tkvB/gDyHr+ZaAUUEyxGVixwDbGuh/BHGKFbI5goZzglq71J/NljKCQ/oaufC
clCj7sptlHSg1DRdxinc98mshRTnUW3rQXvM/C7+PZe9Y5RxqGxURkdCa0Z161Ug4y4fmIrzt9MK
kxdBrFBqStgh0ScJ8imwljJDP7CuqH7AZv8LgdsOwdyvLgeFoYB6u1nbh2Ui0ELvMU+0h8C6knBu
y2773hrMcui8n1hunj70PPkoPEy78+miw3LoSHWUc7HOINiIULKBSv6Sxb/T6J2JUVCw9YiVNIRo
FHM1X67LCaa8WQh21LlHY02OpyVFI81980IrZod/e9SKbY8RKinKeZAfg0dl0CrmKVsI7C/4XySe
Wd4xESrJo6kzsnKBoMyCtfDKwdShy10i5L5v9igT3LGX4FQW25uo2aSILM04UgX1kWLJnnxxX2Zj
burJbawDyXqBf+eVYRYlQWsgacnPA974W0gLF/ueMBEhBIasfU5SNfPC7KrC/MS0J6lASr18u0rv
3GdcULpqXftVdHuengQ9IaAzRivS9kep7y9zx1To7wtZxNDvK7S9W/BBSuEeb9YBNrHdcEPrxCUp
6/3pw7Euprl1DUfl4PpJCmTYzzWUyf1K4W8IKo3fvDVmgPUTg6/NlfERsUGt7qerp012upzU1i+j
3MHUON1BaycMdujCtvu6hsS1RXYlkfkqfDMf5Qd9tgC6+TTOF1kVDB3OmEZSRPe2TGFLwpje6vcz
C3/sqLnv/oc8+yNCdCzTuwTsmBt+rr/EpzG+w5NTRxeV+oMXeUUuenwjN5M/q+bEfGXHJfzqJD3b
k+1tAxhNTtfQA0AeESWI5V6Rkkh6hZMeyKPlgdJKzogKCPKOmtsWjNqX+pKftXQ5aOuouc7CdetE
upXHoJ2nsQ2+UZQR/OfTmuhi6e+WixxUogTGvvQVch7iT1oYqG1TTuZ23YbJt2AbP5Zrlfmk1b2j
C0ECz/ULx6lBph+Qqn05hpfdMHI7rg647/JpYmuVFYoPauIUBlqjkIGaTbuPfSUApJgbJ2dd5Bss
tlDYixIly5JQmMJZ6qbYwayXiMqHfk8iIe6d0liui0RpYR4vd8908SucLVpTsiGnKc2xzlAhLBk2
TpEG0kZnyRPF4TspNhWKWYklOM6yWW8QUHLr1BTUfdA4hdzEwZKUcVr7s7WDK16p2DjCnUj5eAnL
1VA4HXT3nOKUAYk1xHUcPZOyVUcugsvFgzDZHgBCy9VBXeecOLSfT0kgyfscv/o0By/om90BIpCl
VFD5ttkNESMWETPhh2eiTaxfLoCrT3F0NugPpPfxhUt8UDCJe22x2T0R32u5szTVTLFMtfQuGq/W
XEU6wBSyYos7YE5xjREkAiVQ6+6U1o8m31FjgL8ILZbi4Zj16HsXBqu47B68LRX/gP/gT0txryEd
yp+gt/35J+HUIFVfZsW4+nmZudcv7FtuZKomQY1w58fJzwwSqKTOswmiBETK7tS2/MUo/IATNIwa
nvS0+/mRN/zXCS+zuTZfh9Jt+glOY4CHyXl5BM8BNLcEeg3CIk9VgtCYpVVdkWxyns79uy69puMv
IGFYuS4m8wLaM9fiJtILpdS76FUiM5aDhIVLps7A0nKzxQ+ZgDD46XhP70k/ph4+DRnRW0gQuR/r
cT/T0s0FerkNF7Xzwbh09giL5m2TK6dpQN/r3rg0l1n0EQqJszICKswG3psxGhxZAFsvc2tzUsUy
hNK2oyPC0gGnZgljawG5esP2559GmfIts0oKrLlO3vDq3s6t/b8Fn6wW/QcpTXVP0tqYDBKYVVKf
tYduBIK166E2WqvZ7MNFzIy8looxN673RCYtWHQcGydFCia3XWEvAWBuBlI5jv2dXxV8GekNsP/a
x0VzN8x3Doe95au6v8YI7Umt1NxALBqhZUpcxFKMXDaIHjbj9845nxNlCO6vTFVZhWfzVVRO5rk6
2c8j0nf2PKF4dRjo2Y64o1pOoNv0x9JDj0zvICQ1EIjy06784oCi5dQv1b0FtGAwELnI5NcRHGVc
k/6xGhtjkNQpPKMOCvk1LS+sugqqxXAraJUb3vpLs3mcSepi4BCjF1wfG+Ddm21MT+2RWJhAkAKI
voaZ4Avya0XU/WV9VZy80WyVMXlcOmRib6vLkYbi7XEtYQYY3Fa2PX625RDgtDuEMGZ8ZGWViebA
IecL4zbHgRyD1R82yzHpuTwyo7TN8cJ8vj6r9n+ZSKLAKACum/x/3bwl9Yeuke4BWp1xudfqO58u
flx0m/CRYhrdhhWCus4TQxs9DF80jzTlAgIG3rqJzI44/hiqhOE4KFg+CBYMxbwjCOLD25MugqlX
SoSkmyXZ6L4Njt9T0YuMuIt/fPhYWFHOzjHKMlwnerDf2xJ+CXdM7HTNgr0F87Wd+LOoXv4FYHDA
8xwuoAsqy9jxjlIHjtsVcssnT0e+8eFJbL5N7tfmT8lDyqUftCvPMCi+dLUz/483hoCfkTgJ0FRD
5N0YMK4SUrW7fLj7TB4MzYOocj3oYLtFfDPx3b0JX1grMjEiKmF/ZbE8u6G1oKsH51R262mUT21f
BA18kG4wGcdKYGpfAyVm5KGlw6OwFo+g9mMlI59TI1xBL8l1vnIjXMuQK4/e/Df9lbC9zbVbLUU2
OvN5k8kx/W0RulryJIXesjmSa+RGjj3F7gXN0wbaFgUilISpl69r4rYUMd5vLNq+pd3pNTDYkcMN
DOI0vonsMw+BOeho+5XvrzrCIE6hCTPiKnzCdhbJZHAAiKqY/ACprSxs+vDR/TNjwlV+Fysn40D/
9KnlwmdBEkCa74Hbc7GYs0lk0CAeL4OQaKtd2WQGQGyCAQq/zWU0zQS98AYj7bsDEtnVtb510LvB
8/Xdta7+xdX/vr0VQpxMqgmuece6vSatheh4TnqAdC1HcU9GrUY++gx6L+3B0cUor762Yr9Og9G/
HgdvdsBlgq7AdRolvmAapb3CdjhqSWJvEmnA6T30K/AG07afDLBZ6NYUZtFYbB+QpXr9npkC7iT1
p3LPkRZicXwti6n5dyifr6MVhvfiuJ2f0eUq5PIusuH3SDFbhfl1IRWnO590bXesHj5zc22D55Dc
3Q4Og4LW/nEMnANeBr/CtVtU4gWRPAqN0WfUm+j1RE/rG6MrBvtqIj14p93WVCgo1yotzCoPKYWI
fv9o88nsq5onj2wuSfDYU0JgNLW9wJseJsTdXCZKv/RjLXe/Ggrn8oy57uwkMHhjPIMr0iHMfSOu
AR9PZjGWNIyCMHw7yhENKsmCP9Ft4XQfYqrVy1t1ogefSG3NtifCZK1UNJefmsE4+p8yA4K/iWOs
eP3TC5E4yWqbUH3TPxJyiccN0o+O0L9wrsDj3gq2MEAasCpqk7BDXrK9LMf1EYfEuOMdIEBUv82G
4psYjvnygwa0fiUd1KMmHtHiWbH9e74FcqHEGIbaS4HB5OciAOzicWub17lZeJEqvXuuPjLfocva
A4vkuaV//r8YbInAUvgnF6C3zkGHZ5qkCZXZs/q6d4j3gJebDeGBuj34BMggPH8fLLBdjLKiD8Vb
WgdQ4z8V83UbEc1CMqcr4sNsUEfeLpEFai28ve79G2I2UoOIYg0DJf3W3zREPHnWNBXaGzJkC7kq
SHiVKTrWvKqn0YXMg+Z1nbgkVYNKfKOW9iPMfO4oLhGs+NhJMybcxdSLXIPMinhFX1AbmGQQCVxw
lNoKiOcLnbERq1o7zRL10YH9FEKTxybFuVyms6g7AKCL4+YGvkCrwihoohrJusprgV6ElXmA8WYl
7WuJ8QlQWBvXhez0Ur5CwSuYft6hZgHEYVm64/2EOGaMWmMXS0mCuWSTpOeiQMrvPmxj7FmoleUN
Ph2klwNz4a+a/lm+wQCAF8TCmlwDpX7A2Jh+M0rJRxKOgoX23lGj4R55GQd8O7KaWwiOgj+rQPyz
J0l6tzUOnEyaWR2Th+petABTOJvjtdvqDZYT5pyBwlJW+voXHyYHCvD76X7N3yYthfeSnpFi3twi
u9oNVH7+J4lN0EPqZ+2OyxF5yzewPkurQaxkwJ4h/gKoy+vVK32Z4KFGBx2quXw2iYP1Q+LjvQ7c
iayVIrOPv4fbp7QH9LMmNVaLrV9axE4VD+UQhmpqTJvX9mmiNnlFbHiVVzXJV0v73bSLXrCK6Tql
Y4yA+J6Mwpg7jxiXB+ktV207vdw8t/R7PVdFyTFQRKotR8pDycgbuwxQR138xj32+g5N2+va+5XO
ysyltL1WkUiEUDPNQAksNB5oqp2qKGYO/Z/BtKvU5YB5IA6krIHpAU+QyMLY+aH57gGw948vvQz0
DUcEachoS1FjRVMNRZCeNfZYRHl1+4GgPMefUC1sf1laRArmkNXdECNeGZdf+f3MY0NTvHdIewj8
sbOQzr44aMMQgXV55J0/GGHggYxXRdLhKKW3FrHjwM8vVqSYvZ1pnruaGPP686AnuUjF0QL2HIw6
kFUI7uUiPpA8uaiduzNwI1AmiYpWmJhDQsuBXfSCmwQ3UBmop/vYU7mcAEvAH61QPwB3KLPmlxlw
w/MJuGkXjA+3b6nQtZFnglhWDhs3hh2qsDMRi/V0YfkUYO2M4ZoJ+JD9MCLugPkhi9w734RFcp+F
h8HKDKKYQ5DVz7gWeJ1ZD+NgeKGcP7wyKfOeSXLbKAG4K1EuPms+vwi9G7mwmjIxHbz7idAj13RV
e3c7l31qppUslv+Gd3EAWS7SDlLw8Ln98ylbqxDqbY29xmcYkSEP9MB4fcvxKszcLl4+paCJUnvC
S6DnLO2bWFBjG1MW8JTt63ByyA2HylTZ/3B0xCVI7mUo8WHYhGEFex/U4Q0QRHVodSMhsKF8lhuH
+WFMkPAtlHZzoWRAwHmojXuKvBMbK3duL5OytBrwXiQm41hTO158K1QY+JHyR0WpWnz0w/Hxfn+B
wPoiqevQ/kddiNugAMeXpGNFWHxwxOxU4ee9qhNBI6EJxsLS9HKWRXlF9tAzJ3KfieVVg7wNvX3P
dxbPrpKLIkyzGnSu+8j/gDKk1s4lfn/u5rIdogeLCYDnrr3XSWpPUIY7eduX4zeOp1smFgpmR9iS
M9wHgWw+mObi2FxPn0IHnyRaYP9iwU68Mt0/RwhwwZWqRQwObTTvBvBKvl7TGHD6xZx+a7gCCqoD
Zm9pezAXY8bD8PqX/VhuJeEf5M4sN8M4UY3fgTwodefQOaXWPPRgK51X4TFYTGlETLI2fPbhTjl4
ikqN3ALrrCSLsgrLRqJ1RrChkic4YW47kt8bvTPdN+jqrqc4n2AMIAqa1ggncm2WjN+0Tpu4Y7Lq
b15EfVRc/83OxDLBeYdacmRKivyML1u/TWzGxKB1W54TWqYw7zXld9dkhaP454g34+K3lx2Tcbc1
JVfgU5MamyOgTRDOcx+qn37AyKzoooaLZgPM0SFscJz8adRnuCBRLnel+WDzc04jiFs/IUKvSld3
ivEIlKmnshxJL8nPN5ds5vHg/hZhiLMHG4RxyVCK444zgkjckfbOCWX+NxAZ0KoK0+ttIKJCEIpr
Yfx1qD9bh3rzKIsGyYWD8ZZcCkJO6rNqr5bqylIVwONNjVRmmPZE2fhVsqv7RAL6FEhbXxQnoalj
yP+dImldzDVRY80ch3cLZIvg/HDMHvDmPDhcJ3ZMceO75qom7OuO2NLtJIvryQkcV8b1nBjb7EVq
P9m/WjUKuECoJU52mxxarK/Pijdz0whOKXfvFs4Dqex7uPY+z+6IY2C/A1x08gKZFyxdkj07TqFp
6zFb4A05b2DAikgqXLssLOnKh6h52RyiPyi/pwqPVjlA/78P+Qf7h6iYccyIAwG6S1QQA2pNVKuW
jLFjfCzB9xJg1qTws+pgSdANiwpEgYNqnAQHV0xtWOB/7BQj8ovvTtjU6bW65U5rq3oBRc0lK+YX
5xbt//0b1Lw/dhw+cSVyuffVIgDo32MFZ665YH6wzkmEp4oZQ+RJpsKhMWNh4lKhyfGdaaDBLLhw
G/FTwyLh7RVL9tp/2eFWe2pY5fY5OQP6TFzfCjJPHl9uhwRWK0646eDh6w12WPxO/1GEwhZu6/t5
RmWtMBahqFFZay5te+xPQtE7CqPK+ttWYTXiywvb4tgTyTolWe0n56ZGCqpgBdNe/wgPtPwjJlgU
pzmuHJvkQzn1vtseopT5kPRexYgY/VUNdnOAnmh3v61VJ5zgOniuxLF/aodnir0FPJDpCraN9O7Z
mDqeHSnrXmGYD/luYauLAi6r5w8OsaApFt6FznfTk6Pi4Y/WFN5qQqajAHz2SyP5todfxnkxS5iu
NLtT8JJc//pcDq3IZPmp1zKrkE9YdolRZKqn3UjK+QbfvT7A2Axzg8LG6zebEAhqusDK10ITi5fo
n8mQAh8J2SL93RddCIaZwAYeqQAGQZAUnWAha9iMuwhtwPADgdwXWMD8fMtn0CguigxdNEvuDtwh
h8leBnm1DpbxoqUZNswborPgE+C71TyV0g0ee5Z/eg6TNNSzI3DJQEEZvFRf9ZUYxih6hVW5NJDO
PA5MeF+SOU8i2ITBssOKHdcW8UnRs/l0Ap1lbHs9EiM63zk7EBoUqj4lGrBGl7g9TQD8I6VpPQco
EC6NPrFWGN3e2MJDI0DoU922bWK5SY3InWzKcwuNc+UrDeHJprJN3ExPlMDgTpVuujjRJB7828w9
2CyLObWCJNxBbwgdgud5k2GDYAzArC1IvJbPtGkHfxMXg0GRGfsbwqHC7M+K3oYENrPlTAtvQLXB
NUjkATUWJirQe+73zeMfK8Yy4mcfJDlRrc62LlfNWe4U34FraZZXiwHteS74e/iBJMzC0vxNlft/
2c9RBV0D/7asPG7TuukFbWNA4X1VAvF6rpR+WCNeDmQEJJmWn30ztPru1Hcukpt4j8JNZDaYcV64
/+CoD5xRvHaqrmVmofwhmM5lKCTQgiFYVbz/W3vSjWUhfr0ylxQwq1qLsb1M9BFQt/qORYdN3SyG
Y3NLNu2kHG9q7AvvSp5ZDHbLObQXv298GEuU3u6qv7UmecSZpjKVBAP1VKv1a8NWTElOWIQLLHPT
E2Wo74SN7TMocrIYHss1IN0Xfr4c2T6TpW3BeLTi5lhvqM+1E9RdzsZ+O+U+iOj3yzC4nGAi2Mzq
m632HMahtXcKA8pu1xyuHo5jG0mAmN5HEYopx39j2FiJnzPu6sX6OqU/wxtJDjwU2xboMA7W7T1A
MmBJGmm5+SHCYNXCiDSvFLJWWusyYz/hjLF3mrVt2MS4mFIxPIKF5/28qgbcOYNkuJg1Cr4AFWud
QzaD4siO4JdLS3zzsRHPT18ia/F+qIAZGnkE5FsA9A4K9/EdGasaUUuGh/sD3dkmnWoAxSntPSQU
L7/X1QN8yDLFKpSQ8jG16ArmXTjGP79y6VQMRf4mk1Jn39vtYfKpDTArSiL37AxrtsdZq52awsmq
EEqARSQ9W3DPtqYu0ELneP15jBePUbo6ZkZ5zy77IyDSWLxvh0V2A52g/RqvHMIMtiWe9J4JA7D1
UJvo60meIMTILx3URfjGXRx8u5nO32wtX1qlqmBgYk7HJktbBLSKjXyGuNJnkkqZDL88XDtCiIBY
Ed8pi5szkc6PcNbdU6T5pB2qvig0K4/cf4U/R0SealtjQAc5i1sZkf3IOuY39F+kRIWD5B3G/Mx1
tP1egVFcVJ2Njb3HOYi5EJpt8RGu8+B2v0rH4IR9IVme5bD6IvK6xB+cmLlCTL8YD8v5QtO/INNw
rB0ruuEXO1jDiIzo2TFUlaAraVLf7RZWmLicpHpia/sUz1RfmznVNUVcIvcibAoBBIVEWR5dn0cg
ehjglWWKcoSOi7yiPJvbpip1sqKNB0TMutYFbuHBR9TL/gtgurcMScr2aLaVTBWZKfBRI5FWH7fQ
//nWZR+npaDWlHRzMdZn90bx00RGc8uSq/Y4371paH9hBRmmsZv2mUt3Pn5kF4cmjxOV2zvWi9/O
78OC2hKBX/5i3Jyvj9/IBOmmr0DmGQo/zg1D/RFLzRvhDa925RlwKCuPPT0Jc3LTx8D7CL+cGXNI
2E0aKEqB2B3rAO7+kA04ZHcWmgJeplG4AkC0Lbf4cxQfbR6NsFDsNdylKQytDuuKcgDW92Q4ciHj
AMQqNKxHRe3DpIPhkwShOmiE9hqvmn6Z2buGLJhaBsKY9AonGGaA9FgzzoXdA2e66NHA71SNE2Me
Sol+//OV6Et6iljcDOscRRjza8KXmwWpE0wG+BQSxvlX9FGjynhRiFYpgMh9LUbMusxsFMYfWpHR
6p7N84luemGyOxbdWDTENqgezLsHSarWgArJDLOkHQIIpzWbihWlAg4h/XyYHIq0VjUYIxcGzBwc
7JpWqXl3MDeSb/zlsDY3mJicvA4MlTu3o78RKDAnRbHz+gOPKE1lVB6jPla7XZq9NbaT/uAAJnCt
nmAVwtWVsd7a8en71OUXbC6kaTI8l/ebvr6IZOVSaiomsN5WyCRCACHxYw8p/OOOe066BsgKYS0A
izasojNkWu4P3gmwRnioQnHyZcQqz0NMvjVshODZaGrkcKgJv1f/Phn4Ya5If6i9TQ12gcxtp53A
ufWIWtZ5IH0Cmvfl6mEB2px2GJ2UPO4xFwMaqdYwz6SnRGljvPdWZieeIq5WpbXlE65T3EHPR35D
yu62wHimO2lkbCgETimE7mgndivmHP1wXYf+X5GjpmFJ60tV7h2BdP/eumVEzBksP0qvbnVQ7dBA
RFbJGbY4ZRWxPaeEUgmuniov35E/bmpGhgwQ0Scut8GFGUgP6P7eg823DJPN2poBrrKpyITnrMNN
+PbnqYGdirlsWdLxZhvBnW131Cvh9v9+QQgGL6TxHp7fKj0VA83orZHVJuN4gdcNFEbBnQO7Rq35
NbBWyFhfkAAHb31bytYk6DFyT/IZ4EKyAP6Z1rv2WixbhP+wwOtHQEGMPaJvgjRjzNk6axvYhrv+
ADsJS14p8JpOG64PDOe+1glH0MVu1ZoAUUXngpUxH+xgWjVjftclU9/CZpMQtUt13fo6a6uerhpi
dnhS29mgGErOzn/BtEA2ftWakR4IzvB2uI29OeTwrulOJDqm/SjUfOjvJNxV5PUuK+BGc83R++8y
Cb/V3KFy89DNFTUfGG6a5GHkTuQuXEv58uuI6KubOHLyhoGm9H4hCOANPj6c6HtCApbsGBlNsU27
iw9sIOkck/ps2v0fxPnpWEIcHhjxLorj5I2rGogupO3Hx0W5N/w+wKHCH4QkWYgzCfvo3Jl8oSNf
0AZ9aSPQ5BqbZ0jMDN8LtiSZjDBB2Dfypteok/b227MOfBPUWrdTXXA/3b/ZavNiL0x67WfR+lQZ
2LUr8dEeFbLRkVPxFCkpBCEMvtz+7aFtkroStfAAI2VDccBbuTEgkzrubVOgkY8uXH69RU7IzEKA
p2mXUlsNkoIm5qkuQ+ViUxtojNWxS0ui8NKnEvWpz/jfwap8Ineev/O0SSYnlJ76T6byS7QuH1H3
wVktOZvoKEdh3aERZoCwd7uePhgb2w0Niawnai6e4lEZAdxoi2fwRWz+OG/PWx0sUm65MEteg2rr
K8F8rS8nM31I4pD32QNv9PZFtKlLnXjEISoshyXQFBv1MAmrM2t7xaCIny8w25kL0arb7TjfRYl+
ivOBAbWD0lOQzK5Q2BPLtNlZYljL0+0zLKn9VwTF6u7oSNLz7D4aRjpm1yP+ifQzG0dtDEQkHmRi
ekd6zj9iz95j8UjH+N14JlCEtc6WBgEFBu83ZnGFioKhlJ3CzZeDrXRWNVLmuIOrGllIHMON9QDH
UnWiK6tTlhfdLleDf3eARNZABedhHWgchVMfR8/V22A2y8FL+bcjdRNtRN0aw8Nn7SdsbFYbsg6H
cFBdFX9XWP9d37PVtuX17jn6+DXjemb3dUf7OEruOaID5OezLgd8luR+SMeCl5kORrT0EwgBk1Ki
VIdfOQ35rXkP1SVHqnGZVg3DDeC5+ImYRI0CCCVc+cHHn33nXCUUmlv8kgOny8sy3W5Iu0tll9ij
+DcckgGrrDBidpMvFIzvNptjAG/DgINn6Y6UuuC/J5y40Ghvctpvna6XDly9Ygo7Kz+qYiGDH7+h
aQ7zkRC70xF/aPI3wNX4FluYRSlTXsYHkjxSyT2/P0f5U1VvbYEL8qhYS9243TL1koQ4WUSWVIh6
CFCaTVAMGIOfOWoh9UVCNh5v1Z1bV9vmN+Fi/JkIOF0EnGqIqtaAfBCIb/NEniAqdZF0Kz6E3or0
soXow9LysvNgsuAumwfJK99XAecuXgkyxteb/8YDF6UGxAjg/+Dn62q6snhYMftco02Xsdyc8cot
Yb264ocwvzDrJLpK8ImEmTpo8PNKo7+/bSdM8pE/fjFAsvoJ69ydFfvg3B6NJ/Br532y3bp53CXd
3qADSyrf/oo5yM5MBfiSkDSdJ85KnW5UhhK1Jmps1BeCsf3uH5CbNbBe2ZhFKYIqBldj5EfHEaTz
tIkKAgu/rSuz0yIBC7BwQytwHMu1IAUtjXk71/kYOHSKVNFkt8CtBc9rzcjKUlHeMFgZZtvhP+s9
u0bEb50sDhWRTKKr+8kiXlVlPZCfvO8UA5l/f7rL45ZbW6tTYfqBD15vOBFMtyd2gCB3pgDi32cS
IJtjwGgNo6Ia6z0ZFwBIxKKdkIWT5jKY3TjK906woJc9seNHVfQPSFehywjpQ03RTNSZKO+0c+Wz
xzF4b6CGRkGHSc5dTRrUswZUv6B0KtWGjYtk0PwEVmBPHjLigmDEAbiVDc9up+y/dbtl2DJHaSdK
SaNeLuA3ySphvuhDLn5sW3/2F//nPKrXxOcw3Pz9nAKLTm1n9y5VzHFofIvkZ2aUcSkjEuslbd6v
R33Yk2tGHtVDEK29GWyBpOOrmBdIDZbtYhiG6m8yvt8Q14fyMC1JuFkvQvpotUPdL69zEnuGn9Tx
8u+8dEiP1/XJx3K5krxc9K7yoMQ0aRUjYEuW9CE8wAzU1ZNNWCrilpSB+2ITRoHJjTirAbdXGCLX
eEMeyckv9VZscJRjUNWQnxniRt4xkOYKINUpusZToPzlEuo0hoiyE2Xm10Fkat9laH1WpRIYvWtO
OVKAVs3BVJwIMr68/GkghG3q5Z+uiPJmGiNmY7eYQY/ImbhKpDNRcFiRz80V8WX1qfYRiL+LpLwI
8F4YFT65wQXb106RV+vgAWmYxKlSSUVHNTinYSqUoeBNyz5BBtHN8S40n+YR2Uz9GCcuUFbIXAVd
BinZ25SDJNZOaVlxxkEef3k1PTZxChLVUZSATkyKOy5dYExVRNW24J0WdjiLLblOnkqZ9SR3aHX2
B7r2Xd06IjVQIaiaU2OGsI1yLOZ04i/mDw3S91ZzpSIw9UWMfL6rXTUjKu64LfkPUOWDnxljDP7E
VM9SpGE+NZHOdpWVTkMzc1Huc3LFXDTs5AOQdC3j867ZoCUc933n/bKNPgMN7BLl74UZpUGBPGDy
PH1iNwZX+U8zc1g53llQbEnC4k4Bxwc/q+CJze/ZwIORQ1lkc0I2dD8kZ0DTIa13jkd0QynrDcmD
1RlMR9G6tT0RU02Jj9aXBpOJTTOZ5G9nYIeoaroNMPnUVUxsEH364pBHFbME9zV36UJ+GuplcsqB
h0Kwrwt95w+cVDu7MV/ZBmxgY4weck2ohpPTvev6hLbw/Dt2sFxPlC9ewVcbzUQJuL5ttxW7FNpg
sfNGmq2QyndDNmwNrFJYQcE2C9plX3mDS5eBeCgqbQ4dTqHw7e3TGY3v/FugEyB7IfPyNOri2eDb
Uwi7fP2mrxP1/tOYwlm9VXPfXc8rZJwvJ7wFXJoysMm9N2/Pje4C36RsgkiY4kt3RdQKC6wORJ4N
T+atdeTAnJOVQQjv9IfIVUzlmCGFFvHJJOVbeZo7NKKJ5Hyf8gXKIOWHtdO2sJftEadjwBwdFYQc
NE5hjAVDWzTRtUGzNuUnB+MgCBoLueETxnW9kgfIALqLm0B6TKP01JCb+SFoGBeKfudv+x1yghJm
coI/vT4tuBNTZO+wcJ/6xGtC+MGdiMX448K2+WnwFgP7ka+Oi7GJiAcNNsFnE1ds6OpW69i334G/
9MQv3Cj85QA1nMaHV6XWVtHn7DGjEqo9nhKInchyvGMIwtHZqvy5GoZYA2EpZL0uVXzlh9eBP3qq
ltDPYrn8jaH1ivvOAapc9+fNrZ3cTErsjJcoJHcCwzxNgVmqzmgxxDH8jEtLRKo32q/hxboULrvD
kMF8SoCGmH5rMQiVh07C8ikCT8gyGsI+De/GB9HNyZrUQ6FDKnsC25ofhMnx1g0C8gZbASsx6ZwB
C1LOQL2MyavLbuHBm28u75ausBwkznTAeb50XSQadWTeyZTAa5CvDJ/rhTTqbd5KwTM6Hn/QMeWZ
gr+4n/FOgf+SwFkxMp+fL3taUnQMWKi+vvkH25CEAlSeNbcXAY18DPVxxqX/2IicxE4ylJWzwemr
+81DBGQmmgDclMOLHcEGm9mjNMWSU92xEC0MOqrHBC46G3i4NDberDRiIc20sUV8gaos2MZeiES7
/tX11Hz+Atf4GmD9lDDQGNspu/WPcPhCIIV+ie3vG/U2bPkilNvdEXBjDyT2tD0b4yN+BRPDeJ73
eYLUCYeyHAeWEVzxjejnvDuHFvw+00B69rMU4q9VxMmharu8li4Y/C6kZNf4lXYES+sdXHDk9l3D
Km7pWfPAu4od/rQ9VTiPsJFGEzSQoUwd/iKX3okj49F0hkIsov8PRsrniK1M5Xxuj0X044D4aVDE
iy5qpT6yDS0KQ6PFPk91AYRE6ecNg+lRIiu850JQzPh3CS6gAb/M6i+KqtkIeYYvYEBPP9SMWO3o
XS5J6hV8w+SGCqHuuE7AvkW6wPZTIBjLPLVmiR89JZukE09+BBVdC6+UFbvLp+637zIfIF4yGK4z
nRq8yYFdMD3V6nEWjKPwEgdWsGRW4jC2OvYDPjsSzbobl4brjQZ0mDQShslfrnFzT8QIslUL+2uy
zD24W8eb2zmyPWIsT4V246qrt11fpiHG8IeueswD/D7ywDAlcnVwiy43vdtlFutDT/FxNpg/OUuP
p1MZVEDNVUc78AVcRCUEsTZWt4zmv0CL2T8b3DOz3ZrteZZKX+qK6rA+xR+3UL4e6d6Xe7PUG6L8
1yeWF2BKtY9wpNE5TTZNhzexwt3NFmtrbK66VdFMLNlzpJf0ch8Ln6o6kMCvdW/AhyPYwXHBTXcq
EDyKvlBVOovliElMXkGwkM3IilRW/jRHhXSSwRA4ZqECttV6D9MvHMnur/4OiRYk3MHd8DPaoN6t
XwWri0t2C2I663o9vPd/I8xKNJpWSOqJMxInJr5z33QZRUaRaYGYTePuXtVFRQhkqE2Rwa4DemN9
1Y6cBvp0MmhrxWc4zgbNbmOz2H3XnA2zqLeBt3DRl3BLcKHsceSa7E6G71bkqkqIWTPqQZ+jlvzT
VSCIgtyPOdOzKCQt+k7mMJFwoA1V5/pGT83Rc5+THQ1fjB2eMpkIHxxJ546FbyJ3rsv7gZphyZQq
thwk3NtSun1taWtqxGjS6Rmz7ZEtqXyWXf9z/vUaNGQ9yjjxkD0FhKVOa/UY228F5V8qNJr7Jawp
qjoHXAmhCEpkYEer7A9cwYvPKGyNMObP6twnIkPsecCbFOyStOHtDF6Z2QAV8zincN/QhGgHp3Cs
K6GNigcykNmqBfoj8LbzIlx9uIr25YCMhaRcWQhaZrIzhsn/G3kYVucsKMK/VQfHPK2LSLD8Db2t
LXMBJwSRdLLWSAkNVhlqkNCDg3UjeQPl3ST6Du7a6BdBwkHukQFFQ8LY5kvc294OfG+rTLZcl6Hg
agWINhRGcWVO3EE0knTiGDNoXsSAJJ3K/fJUuOU/t53crUUk414KbGuBbxL1cc8gLk+cvFXjXHug
vpRmfayrV7COB3RrnKgx9hQjZqYoYhW+JZCXOv1POxzNYaVAJ01F9QJTOpPPzidSQX21pbUp77RQ
Q03OnnaNjwA5j5AEnz+NKToeAJ2H7B9+AI/HZX/vKKZbHKGgiLaXNBE27kWUuSYQKdqHl8ffVxA8
IL3EZieUTnXvZyb2Z8WbbVlzToPBfc8E3DTsBIrlW1E5kUPfOiJtVjwerPelOZgowFkLqCuq1sv7
ChgN4BOgShXINte594hd1B0iUNNo9X2cNfhXfhiDlWJ53pzF35bonNEDOw+e6XNVkY3kZPh7Vzrn
rN7E39ifVexd+m+Emc0Ke1qkhRzggB7j3IE4j/RXcWWaOBbMOiiQlxSQekTfGNuYhmVkBZdOUaLz
TGtWiJxN820p8dWJ0jme0g6m/j7qehnr2oA0AuBnRGsGVYqyDxXGRC/8DuS3Uk3GTx/N37fR9ZE+
3idBF79Jc4N9P6vp0tz7IF1oFfs+AZzZU8iZfkcPg0ZijxLeyD6RdlN3wCiRHoT/J6TWEyRee8ky
pjfz+XtDjc9fQau8/PkA0FpiPkyD3AAKUEGo61XC+5ys+NIH6m0IGQ+eBY3zjcF8wnkVF/M/AP2Z
1h6Pgk6W7tweDvaU6hSLuR8EbX3mvZmeDzlnTxJuCHN+tHas2I9cYKWFFxICtGwIjY1l0zm2MBTi
tUTwF6n+CngTcm73STw+k28Q5PreyTpWkwnh9kWHnew3LOIMd1BcKdWnWwDNZ3g/D8vqNokdI9wP
DsQSCIfPwSCheNCYihhUQVxQxe3zelxWL59FwDXlnAzvgYG+Am1pQfGqxkabEGRmgZHfC8iFaAAa
JEha1NamP6rksepO+orMBF2lo2a4vpV9HQJbwhLVrZWr+yp6ZFVb/cB5JZfxvKiJbZ2VxzdqHBl+
K8HRW4JhfalwspoAILxDSr+Cw8qrBuw4bxCwLpwcw3leS91vLrTHG24VRFfE2Vw6w/6ndVieIfHo
sQS1CF55ImJfn2JVPb5ywWl0Ti7qzbLob0nHx9LbUKP7pPnIPq6u+NBQqcems3gaOd9whGZGy+Q8
AJDTOicGiP5m49DXGU4uXe1woYvTtuvBbMDeg12PjP9Htw7VS9Q8Vxm9oJkxAuCu6Fh2SyYOdtL5
zj0NbGz/cI7yEUfsEEseh7sz5t6ofxEBPZ0mfgvztVYKbr4d50OzZHj+b6lFMcVLh7VCFGP4ophV
Nw1JF+eWiOGPuIYLal4GfUZTW2nHBvQh/5r2F0tzCtBJn71JtdUr9xkQqU0tzwYbsp/dpu5l9jRd
OjLOKqGdTMoJiVkfaqSD35ElIYigk/9DhHQThvXVQG6XG+Dr5F3zJ6CHxtgoZLzrgRvMgRmOfWO5
r7+IsJG65YQXMl0A+NuSd3R1+ZK1cMvksjuB5gfqK/Ldnm11IQqc5TK98cEL5RrjcDma0TDJn1LL
repM99a27EwgVTMnnWm/FgEP+4EZqwjB4ThD4rXFCjH4FmyxwnK+gejsDh63oZ5SmV7z3IZfsEg9
WyB0yOSIP8I6uJ3CEVhdtUIbJ/uPLMdd24hsGxnB6S+6DqG9iMzqIocJYoPYpdkOmYBgFxydGYmS
QUl2AsYsrPmfywZ5NMm7ENvNEd1aKUMoD+XsDtZl4eDsOiTV9SM/hrSrlweGHU+37TFK+3hGSG+9
fhwBruQbfdLeNyGoi03BAWPyxTI5IHSgqkyqpnVU6a4hiZcJaF3w67C++GDTcWRy0GzEJUhPy2Nr
viZV3Vqvmw0uYI/CpNriif+Ro/67dqUyerTt/wOphnDlwdnwVJzq9TpyjSTf0zuqXOidazwD7dXc
nv9/lv0RiMc3hbMPd7ADxWBb2O37B9UaC9kijGVWazEHbv3EALJUGl3Xsp6RKT4fIy4tbXdznZnB
41TltUJDau9EgDr4RmlSw1ojENFIskZBw5l3wi5UNaDMMj87iRutHWb/ybpLvZcx5x5TLPBtnuX2
kVyMIPClfPPQAn4Sjm1hP1qLYYtUcc7B1Pexw3QnJ7B21JAJOj0gUuVxa8J+JPrmOtn2dZLDkhMK
961sXOWNGaJP2/n97lBOtuy2hRKBcAYE4Eet/fdCrohThvBx9UZlWkKJwcoTepNX5gL8VnPXHbMo
x3LxTmlNzuQbcOXl4lZQE3DqOzoDRb8+MTVZF2GYwTyr14lej42lSEBJ1H9Otoaji0TNe/f6lGf9
wjvfDOgykrnMO6bdS/LAUR03tLi0StdbSjl1piXTwktDq1IxuM8taGwZXEWVgTyZxroD6ID6R5NR
vTXvy8MDMCTxMIfXgjiHH1PpIIBt2SnQ9GeSHLlFgZtX2I0yz7bdDkr40FXlfLh5vrluWtkLEteQ
kUCdy8OFay+XJ3VpQMzq88nk/l4MzvXJeurdzFIPy2jU2CgInLvvmsQ4eQe6skdryL3MCw6uwJWY
YdVNacxSUm6oiKlvdxN6FSskEVkZxbTBGnqvdvW7EiFmg4VFULLoxh6IDPCMAzO4UwH9Om1omUIh
QORMbqG7UcH+hZqff8Iez9hkdrFOybHtvbvmkOz71oVk+2vU7BOGT/RwJlvqt6LsUvBjAT54YSYy
v8E074wgS3xrQOghg3E0yaYGb/cpFq/WW2+g4zsBAhKYlKCTR795zvKg202Z1f6kQp52+HlBcZ84
YWBlEfor5JWYwXgZSNL2nJo/YjpFqmv1nam5hWGI+NLANEKFxt8Ye8l5oz4mzGODjvdPM23R0TeU
TsVcPZUgIV6jiZv/3C0yS0VC1sit5ssZRA3rdSf/uJGZrBSP3STUcojZuFfvuWPrRUR/LSOTqbhv
W+blOOvnG2BY5NxGV6nWrniYTdVqvLJZHjGNX0+mog95WDBoSXlq9j1xOHeNCFJ9v9PcGEOonj44
AXjPN2IcYz7OAVb4v1XccoYb6BGaLw4tZGw7kaIBW0samwebiqBSn3GCT60Y5QzDqgcpbvSmHJ50
BHw2diTBPJs6DmiTpH1bvCgwhj8b/HLZFbBQdofWLN3JWO9CGv0PzDtQavZH8Xhse8I4Vuhl3nmT
E2USqJxAeCUrAdLPyu4kVY2RxYBTewjoIOeu8lR8p5y4HLLco2FgxrunIBShf3J+iIin1TLeUOuQ
Z6FXv9eXXqyO57VNWj/s689LtHAbq8r+RfH8A8JDyzKn7MfjjHMU5g3VAA5yaxK2HHanr8zCl1/m
REyTkFkm0FDOZ4vV48aaD+Hu6Itmgbw6fawknl4hKz2YnXY13L8atiDQPkA5icsHPD5g0ufToGpn
+4PLG/6gLaDf6lGVMRDlQvYnHyMqsXTce+iJfEgmBRa500+M55x/CqiekwSfPRQ1aeR8MNOOc+1U
m0NBsXSpQOcxo6nZzNImdlDeH7vs+EzGqrhPF0CvsBkFUbx90UNsgmd4/seDfXx28zNIZZTof3IS
5ym5V5P0W6Y4nRTf8W7VKLrHj/6VbQ4LwjW3ARz4d3Af0zM+llKFGU5KTS/itrM/UK/6V2MByLqA
obDOB2jws8jwf7uDZjhQH/pROV8ygjD5xxDpM9bO8nrQ1uENi1c68L4m8dZ+UwmnsV270Coy6pgm
mai0PPlOcYUMphiZQ8dc+Or2c48dKuso9Izqf0sorPEm7NjLaimaCYTabAT/aop5C+tooJiz0rQb
I0l4VyzbheJLgcQtoVtfkkzO0IQWKr+pOc43m361xjw2fwlqro2KBm0887TqkpDz/xdi97eygs0a
FEmz97yQggom/HvyRQlxocz6ziIJwhRiE4WJiMuWXqOPQvQ/yXCqMIcByemcjVGC/ARl6oM2hvv1
jNHPrpIc21JPrbll5An8+n9QFmIQhY44eNFJcH4mKcFDnTCzPn5t4VIbqPUq+IqwcsZU8eaBle3+
d3bqqlxdQIFcSY6kqWLj+/THWjKvgRDoAzUp2wM5iG4pSghuHYHzkXVEQaLayhpXxlcVzaHqwUUC
4z0Qf+srh9TPJWi7Be4zSQhWsvh/zxzJf+HK3n2FjMbbNw8nhX3xsjVCXyXvOfod0c/JAdKQR2gZ
FdL0phrYJzhK0RbseN+I562yrZxYDqEDEqjWjDBrYg2VSJUtbj73/f3lWze0xuh0ECf6SqCN+nT3
iPfkPF0fNS3SuL+WTgb8rYP6u8FA46FsJTvxvBB0nexn2lvXFKuzuzYPKx2wrj26RGKvk/RxknAG
y3sqkJKHeFIEG9GkUQRNjtF9yK+/BrtKLT9UOLIQK0ZCkKPcTTpGDvn0v1AvH9LoOacTwDW2OwPw
Gh+A9lowAvuibHULLH/6AyaiUh+jSSHxlUr3ywoLHZA7NS1FtfKRrn8MZMLaI/9ywB4wXzIxzp4S
OAx5FsyY75CgDxFYTfonKWsm8zYV2scqy7E/6DSgo35NTNUV5M8vQ/0i/6NBVGShZPb2RggqMFfO
VM+/xIVUS4tcYb4dLpvMP7BuCIW/7MOFOHATjQHlDQQ1O0o8sATCo8fQRhYeLZ29/V7UKwi+5PpR
tCE7v7XNWav6G/Bx35dvnmSZwQQcH4J+LgiJdhdDdfkaJOdA43Xv5G6YTWbzNRySM+SJSsVdV/vT
6UYXUSYp4GsXclbHlgkYA+t5NJ9BXXMxoys3wSZaipqvF3GKVY8YiDyKoVIIIYTvO643mSEWITUb
2TUmMzBHXUVFm2T+cFEs+9RveDAiWQBNwfyq+r/8UrgKiv6g81v55Tb16PrDcU+KbLAebS+IASu/
lP0MM/pRRxG8WLTwmXbxWGPa9DwIwZBq9HWIoQl2EMFQDlRn70GKoDUm8feQFrJ6BZkU7u+W1nVK
pZqiWjny6355tnYCb3w6QIxNz5r7pWBh59eBaQoZ43hEE+D5RZC7N23FEYnlVPiX7XNvtmMDqNrX
2oBSDZikyKjn0PpDXxCVemzLwsHE6Ift9Qmlw/ImMO7dkEQwqiFd/DRI375cWATukiRejA/a05Iu
gfDD8hQERrgoGc+XAccmspXLsLjRgiPWU9eufuYTlNm3mC8GrGA2Aq0719jcKT5qDnMouyjU3gBu
W3WMC1U+dYg/g2krmIYEiUkc0EQIOeJGFknlOlQbSOGHpWFUzcBc/jasiAe8VWdSrB3QtjhmciwB
XHW6m547itW1MvGm/ynIW6j/r74K7lM5kmS39wj8cz/cL92fFy0c38y/wqBDVRlG9vDnvl+5Ifjt
5rc+j0GnpriA/vZDfcxCUWKcysMIxDVzh8ZSBycNwFEKeiPcaKrimvPIBhA89LQv6T46N3+NiGr+
4B5RVJ+PBDSNdcpn2G6A1Ml2G0Yxigkz4gTDMy5cdQcWDd+Y9cG/z99hYjLfEZrIoc/JJjxRguej
UYMccDxbRe9X1RYifuqAa4IVSfVFSnnmF06rWVru84XLBFv0F5WtBCemaWkL1SyGJpFiZf8ukBqZ
TQd7sTvF0pk10V5t1uCS1Kfk4+8SlTVo/2J7XHqRfhQ9qa8nnSkaiUG0/mE1Ok7vMcWhgrHOCb/7
J4R0o5Gqd+lOuSiv/4uWXtG6inJ9iosKNpddEzOqsyRCmfzDMUtJu/LjK7hLS+HhRYxOMtPital0
NdIiSSC7Z3ZeRn/qwDDctQWC39jXcAOJ4u474zI1Q07CUKifolbzyWrvxiiMAc/P1baHOx1l8SDr
mdQeb8EGm1JmxzgHEOA7fLNtXX8YQBtnrk3eDrBjy3+kXOmX+6K9PaeNohMyRFkQKhWJVWyPihHO
ZSRw5QuiXbhy5gyu52uLTFb3ZYwFvM1U/khxwJMmYDj3y8bzHN+M+Wn5gk3f2ANE9R5NhnZ/XxDr
dTJQYxv9ppkn3qkLm2YyVZr9JTlfO1y/lEij4W9vf8MfEffUNd0O2F8JX8k5pxn80JqvP8r/URgq
B5F0LD4k7ie3WqY1GvKAAzUAkAHdanPGPzQw0E39rIQqDLgadKXz2dkAlKQqAX80t7J5KiXPnA7F
C65sBsh8al1XvwIvkt7wwlbDP/ZiAhLwxSqk8eLIHqtAFCChXpBBz3qVbTUe0canoXyd2DlYK+Qs
K+E0VStENbq/RsRvDiKTJCSqVU8e7pELwcnAiWNfDwmj+EnuXlLo4YMOy06nmND+rK5gDgOgBUF8
+iIOoXwjMvlUqNYFMCR2aShexgHRTPEsJB/v/cz3TU+xs9pMdjS1RB8GqXc9lEjRtuRZFcD2Jklx
v+cLZ3aa4/h3ItC+fVhPNOCm1+GRVGxRFjVPATuies8JLix8godp1yIXMYjdA1GKF+00FsuwqWAI
8WJWYgDgPnJ+P7m38mOQ2qK5v9zULlrJDhY8E4RbuHNDvro3BnPGJQfTT2THMZhHhLyuVKmh0OKB
T9eD08DjyKSF57xdkhDHd9kGJCUgKsE8hGUa+abLjQD+ipM7ibar7fd8WVTMs8WfG3X5YGd/DyEP
F3GsQnmRZiA4fJN+Y51czOZAl589u0Utg7QY98QC3wf3q4JUc7taHp+ZbT690aDooO41CTzq39QD
5kVwHfzi1TgCKMll+Gp+0X+NznfzfeQO151tj9qNHCfM1UR+y5Rqdm7rFzuM2SA/H3W7EQKqKNr6
idq8dSPIOeHx676irDR+SC9+Jd07DwQpd/vr1OoCpS6gsG3fYbBvuiukDnc8eyLgw0nEDBusQPTw
uvIKDHHXt9HTj7D/ELT003xBprc4K1Dfc/fV3SAU3By9zUlO/F9HguhuKf4uqJ1R9JlbKg1bYVjW
Rzm7SF6IqQPpZRjmJsc6EIFCclQua/CsL2zOoA2YGTc3QXg16lGNjnuHARGsLBEcNQnJZhTwdq1G
23L3sloUbTL5v0ihMd0qPAopbDPg3Ny8DlhpwUACbUZTzMKmcUFG3JUW/oq+wfQ5uzpiyY14FN30
ImpOMY/RBKZ40fk50wPhWLZyIh6zYw6ZXbXJjt+GRuT1YIy+ZgC0xkiKN3ZGMagkH2ue86NsYojK
nOPgshnnqzkp5XFicu6OSCcxGjJDBauwEMgRr7ia+RXzzLplUl9WHEC6YgDjqs8zlVellrBCvOJP
6EM6U8JLQPCw3HeUVE2dngExO64aZdmrSdD+P/rbmyJftCWz5R3uUGniRcs9blhuqkjswzhmiSwZ
yXVa6caWkw1u61ydTF0in+cLTGzTw7+grn6AY25gxOX9Yrh62Qd4xe1ZUxKz29pq5Fv+PLkGe28G
WVXJ1eQNY119r7F96uq1tFm/65z7Gm2yWSZVPHLwccyPsaUhXCPZqYK5USdKownIzwFAGA99e5QY
Hc5pOtjYkQfmqLUTbz5Rw+tJxO8AfAYYJfTvJeJdJHu+BbKSC9N6TsfeDnUBXwcRPHf1xDqTGc1F
Qn61hYxaZhInpxzb80KSm9DYyhuCc3TU6+rl1T5GGSk7ox9Qp+VVpU/e+vcmpXDAX5obHpT2R8Jb
HF73aBSxl34vEsREHQjk30fLYW+acNE8ikxKL5ogBpiVnm/KIVKnyn16/0cJ6waHExU2QbnjdhOx
F25ILMWfRa+u91U70LDtJTkvGPRqE9NuNf+R1LA9ModdLgn54GWXReij/UtImW0mTXNYvLul9sdE
V5SpOfG53MVpB8CL3qWF2qls6kuWpv/Ezs84u0mbB1eP21MGBHrQNrAY9IWTjI0SvJ4zsQ597b9t
Dm3xZkuY1JCHZJk7hQyrXuBcBVdpvQyF/mN8ZIt360bGGInlZCKQbvTnr+0ar332f4B6mwDRWwJT
94dnKFdtHBsXyFnn5U4E00pq5Wd6Ss6P5l8cUUSCmmmac9dRkhzb6BL306JIYk39LK/mn29BG+Ux
+9G0p8KKAOTbxxvuMOxTvFomkNKdUjTF0KHlnO17TvG8P4ZoQeMfi8vnFsu6SbMZgmpMunKKmpgA
d/8nFLnePJGWwxCJJ/TjjrSUb8798yn+WsTXZMo4KAJFmjcSxjecTg43BWPF4yi6RaVIPqxFvxIk
kETyzP3ZEqvrX62ZStqRhIT7mK2c4/+RClVaFkc1sXZxHXas1itil7Z3szaw/wKVlxL/9vm/fXm8
2cPDhAdGYLPdXGI/5rYNe65AGzQbuigeD5EVlmqLayPwCYZxypx9hRVWJ/z2dyhGp+crX2ond0fF
XdVQPFYrVQOidIpNpmkWVRgA4OSbu/eFDz7BhFkS4A5fvZvGle6H/65SyCkHq7QncilkEb2NyjjU
40yFzKrIJ+kHLvaeDzk6ku1DMvbks3e8YYO9VWVb5bRZStPmKgMGsmDYj2vH4zYuc6x1xmUQ5SdN
pNWi8FiKFgmJa5Sm3rXpqr9K5jFghPTJYyFFmdawuZ5gb/FPlfXBl5JKbP87ZxXCQhzHYu5irvdx
Mh6nHOsaZiHK4rMsNzdcgYd1YkjeU7nCqi1HoYr8LZv7T1/SQsukdqBopG034BLaXzoCM9Ip2E83
hVUCpfv8iRfLyVIOmDCZ183UoQKpuEUtkt9Hl874jJ5PW4EWtjj9dB3319a8GMvSkyJtvFLtB3c7
YMbazuf/FpoG1yOKuqerceF7kH3zTzCayz5lhIzKt8sdFW1VpUT0X/PCDSuNOO+zdLjk0GU0jfRS
+tH3ZaBu9yPVZD4IAxZR+6fHqu8WlJkkAWNhUmopejPmTnT9SKblFPARr69elWTQnRApfxUNG6F+
+PsIOg0DRpIlNVd27AiX70B+DyNwSwCa3GtLZmPpnLGxt9kvNQ6GsVe2W5VTzDfrh4kAxta9N9eV
CGiUJjhpZsn52mtANrrbiaIZldoFw5o3G1L8HtUksAV7mUA9r+9noiuk2oxtKKsdG2GdmZgH8Y72
sAXVCy4uIhNdU4eF+CyJr5btMjFE9J0ZA66KhU3oYIRshGyDdpJ7oiDL7yqnRTGerMgZ2bbH42Y8
b/zNoHgouotnS6k4CTn//UGWv+dRIidmSR3+62fdjYMG0AxKjt79U9CZXLxtZd6XnNTWZB3o918J
3Ky+ViQ6l5VsNJKD1GxI2Pimg4+BU0fpImDuFEn30gFpV/xa2fI6bF/2z1j8o+Y6PSmkHCGlFoaa
BO/RB4GEA3M1s1Rl9QmEbJ4fsxtrxnzF+nt7EUTNDnrSBT3o4++tTtS5w1+fv/WbnHz0GrQ1FgbQ
jsQUq4l51NGZsisG/xqwB9ITm+MR4SYfDD7mwLgrsOZG8MqmtYoyR+OC9aSUFRWs+sunIT+yuKHk
T5d0g7fljs6JM8r2rg7nQsIGlvXdSOP4ZOWESEOaAA2awUpnJlo0vYYYYU3rvOVX9+8sF2RuGDFQ
yNsILce08sIse05H2YggQlE848QHt3AoXmDbPlfm/RLXwHfcgQiH+pDop4wLx1WDprHgPZWsCUhK
qPT7A6oUYeEuTVuhczfB3XZoQHrx7R99U9tlrS4Ni2WVWaQrVi8fv+Cg/KAfZlz68BWhGs3d0hev
y7z4tmO9ewaspcWVuienpQ9qx3rhNULHQyYCgJXtZd8LaaiRHoKY3/5BCVD0JfSuAFpoTVhq0SeA
+oyQAx1WfFhopKRmAzORhwayCRcDt6GHabrVEAmebEr5esATh08NIQrx8plFW/iUBuoxyZukoxXg
zuQZ/24PZnrYb79EL5LUfxiQBbo/cdwrIXg9nItGGhBEGOpassuYuuQoK0VcMUvnv7hHHxUbV3lO
rNXOph1eyWO6MAina33Nh0pZuQ4h4pEhsrTHVqYlmISu1yggbharM+FS0037lplPXx4M5lyfKZAL
bftLUe5FCsO7GKalNwPcu6t2QiYPb2JNOK/TMcpmnGKJey1INdBQjlKAIeq4QUe2pKXjtVAGmVN7
8XSmCxRjEqstROFjCnYWMQrdgbvNhAuxiu9FKFb0GmXSiHhCPTrmBqFeo1jTLhsInToUofK+tMRW
O2yFb0G/uFZVtwOMlFvgaTLX1H8yy0b72GTAkUSfruwG2vAaeG+dx0uHrhqlObflEoH2URJCNCGn
sohsWq7znkQR46gzHKiSlcQIvedAD/yy3fkvwGYpCSGEsv3oTntaTlHSYlUfI9pl+qSJywMBWf68
2OXvXah+itq6vKzPK1NWNpq6bSKnMGyDweNnM924DBJxvShCri8oe05qYgHcHsX0pKndbPE5800g
Pc6OgRGTh5YVfXhAvrP7CbRs6c6vEkN5hly5+r9Oz+Z0SSH5/0wJ2se/fUMuhj/e063x+IUYeF8G
q/luDkDjrIG4V/AXKCjIXx99zkq8SzuYbUzvcmPUOVTK0skOvqFgmaZ70HKpwYO8aJi/y9sk/fSl
KsEIryKVltdUVy+27R5YXV9en/IYrZVhqK5bhNoIm+Fu96Tt6Y5GyLrMq3MG9BFMF3eLP2YKbSaJ
F0/yqxPRTbaqjt/9vmOOABKJ9NzEzet4WVgO7SIVK26yRt4aYstEM/efh9A1uwY5ziGGszm+hpE/
PBcKFIHm2M0+9h1BKyAbG3eZxj2f0fi4iTQOMWfTga/g+NhvcuWe/4E8JuqKfOanJ7sgNI8WTc4Z
m1Fa0MqpOYiuKsmF17QN/qHW8Gui+YIzKq0HaD0a+0WSbiybSj7KGsjRtpa08OcvNESvztoRVsbI
oVkkCyKUa0VMbTMplB9J+j1dD1KyVUX3vfKtH5VxhOnpiS25T+GwhSY3SMIVJ/o4DBcA3JAYyQni
MITadxdOeY2eQJGOJMCsawGREeG1uJ9dMZuxlvStDyrHoWERpjeS365BSUBLn77melcPgSL+Jf0o
1cbto5LdYRNuiLeiPj7RJwliBprUn+izRlJP/2BovrVCWSfrTXXtapoE8g1zkAQ04WBOr55OjH/0
p7AI43qvM0MToid9szMNxeDmXQuGdSYn90CTRXCTue+r1w5Dae/MShVagP4zoSqJ22KblqOjWFZ5
kv04WM74Z3jIdEsl0JIOL5020XBEzs3draDiTf4Qc3L9t8tn6lV9L5eJyXE21wuPepVMNi7wyXdi
SaWI1Qdj71Xlj8fDymx9bOWh+prSTovRUdvSwQkz+KqdDIznr1KO4TaS6u70JpGMPUQftwqNMCAU
yvIvVXkmbVBXMqFyVFjQSk3Ky/ciylLYNxA1BT1iSwzOAQIcsY21o74L//12M9X7AlJJTwhLt1RO
h3VY1ahFQNpPwDFnqitWrCJwAjcXRJWqUdoLmhgGSCdSGqMErhmPn2oVIHMHEsSwzrOaSEmHSOlz
HCLmcfaG1XZ5XgluBdjGL2bl3ZBwmnS2H2FjffdZyDbQ7ixz2+V1Bbw5A02F4ZfAEWasbVo1HhkM
Lr2GtR1PdfTaLH3X3bOdy+JWNXjnEgJybFbr6rL1TPw0HmHZRNcUeG3vYHldpQnQQCUTRohEsTqI
kqD7JdpSSzns/aHtUR6QNc0hfgYRY3Y1ErXunMzCqRuEm5MsO31xd9l+86x6XsnoWNg5AeMsibDG
7AkQlOCboEjy4DnElpZgAT/KzGhaNQimKbbW9j6Vk/4k7+T4paOBkThHUDBJfOMbOfoiBayNxUjU
3FMKr49PdTXiW/kPemLt7xDB67W7v14uv0kbiGg+Buq6Fxfug5veXmOtBprmHsY90VLjIchBsyG0
BIh8GKyrUKCiS8UY9n2XI+z1cywQzZDTQE2syL2y1K9Ex5DRt0lwHi9Tt1mXRORUh5QxTctOo+3h
+/FBGCepUfR54g02yzJB0kGqWP+7JQ/s+vcYVW4zjk9wlvu66TB6BaZTGHUmh/qMYzUNV+LEIWDJ
81C/RzBvFu+kqavu+Rmls5FpW4DlVOXBRgv5udliPUgPE65leFY+yjK22FC4ic7YVTQNZ/EbGJNj
Z+HkDYuZoqPrFRC0HZXpKYju8TGrXPcbSjWxCVoY4a1W1MB1T1yzufYT9lHCQb40IFQfs9QnfTn2
ZizjWVFVvdMleLeQ1fbPT695B1YcCqNL8juWIIT1vtwrVhAlon+l+eG/Za93i3m75/o7/mL6AVvF
KQmpVUNj4KahYKZRJ/yrAxsOfKKZWfqK3SEXx7OXDdInOZeEfDkwBeg4TZaErf2C2Ag+8rQ/rzsG
X8wxW3hV2YepIqfzgADd3oIUplSSc7+x8KcUtFWm08eHBwSRrWlhNQhDu7VzuWB5w2HTuYhdjPb+
X9p+TcDDI2n6qsHV5H67NaSH7RihzU5dyx/nsF+QLG+PQqXQ9IUIl9ttYZLiz6eyYjFRiF0vJu9x
zpktcM898vQSJXAGhRParqB2a+LtRImSpQxymV6qZ7+ndfHNV9vr+XEXZam2nELKbvN2a40GXCpK
lTl6UBeZaeerkStyDaabFrI+bifEWFR22Usf+ZBghwMqi3KAlvhEF1X9CrLj8jtz0Tpw3FiNvweY
lB+O4Bh4PDCPq5UbFSk/+4rXtxNf4jaGUjpOFwIHDueJ3F1UiUoE4OQcHBKUyttCDLCURiKtPyx5
QuAJ90+tYukmFNoD1V0dCIS2Ld4RJoN71ST4NQoAnplc6w644GfLykRdC9JVsGdKCRqqUTsha7qf
FzbD4c5zdFqHlziAPENI6a10yoErChbY6SablOzhFdUrOuGFjA+de3rtbmnQWa8StLrCBuyvs4Wm
Z+jb16NCvmk6xgkCtN/w9yfPlJgdpkRHD3NMxWBHp+G8sciHzuq9Xm7So+q+NctdsvO0C+kpB9rC
Uzn2xDycirZY1e41C3puhWiT897gB54rST60C3438W635FmhkjZSnZE9C0rAlZeCs2xjzBHOVpDA
WOzvUv3+QDeCi3saMqGsoJ5T8B83gVOUxNo4LkPBe9B5dxUZG0SYoDkQiD7Kof101tF3egDt8YTH
j4ZqTryiL8xbFtLIn4VzvEOdGcIOfzVh5FpLIZhpKV28bI3GyG5IgzInasQEUNWo2FD5irX0eVFU
Vfp4V9mWX8gvR9WYf2rLXzbbvO3KV3OfV8lXsy0FIfusRzSiFKLJ6cXn/r9FqWNulRvSbNlM3l5a
yji0UhiY8dxlEMr3e490SJmiomEgeTjbekSW1GgLPkd3em0u62TNmxuMWomEJ24B1z7phG7glc0P
jwk8IjOXXc23YrVD9O1989bwMXHEzT1/K//ZWcHwvBaLwzGD2wqXgR4Dv76Sio3IoMAwralUgAnF
fKw6kh4nR2p1HyjkqdeNYNl6o/mpiGfuGu61ld+cle125gN9I7htlLsiQAsQW4xilE67/96/usGO
cmrcCzziK6F/xcWcS5mkAl26bWLP7X4UTQ7tCtQHzak3iIXRHnNY/1U9RTglyjYfDRh1TqbYGbmd
VrU5jVlgBkt5gmnAEbLKPCrdJkvRB+tuFbezWs5jq4ftmWVr2HQXbRO5LJuJnzTE12zcrLYV1QfF
9+VodnyDV2f+rHZ3j3QGHANHU/cuOVIESnMzqOeXpgckk6XuOj/62OxpIlwtWYkpBTsQsRuM+1e6
SyxeGeSkRxz4PBZfi1Rxgdfr66nfOzlHBeLzukl0SMtJL/f69dtkuzFTjplG3LwkQPty6XT6rRfu
PFM5Vgr1TRrCmNrf7qTLpsRcOut4dmwe5RRFqjO9hKDz7PlzPJYvN7TqD5x0SfeqVem0kdHQBMOe
x65W6Xw4NathFz9omQ50E2RCap0LfMa68J6wQhtz090AG2FWsM7Tb68E/ZkYs1+zF6V5lfE1zPt+
TaPibrDLmHY8Iqlnem4XJxNVLltcXcT22p51qq+8YAOJJ1vHK25N3+sE6bYSmqRF8KBbXFB9oaem
xQWA3D58ouoBPqa/aT1871/8xmy/TQfelIc3UwcPrLp/5cR/RPv1zklAJd4XCvToOCU4TjNQ567y
cq6W6BTZnJCsRbhtNknh/rNRmzWsBYOTa78a0GWlzEEG/eYHn+qyHc+cmsxK2P/DK3wzoxJWUPpj
luK6lAHnl3ofymkVmEfSFPYM0D5k4eZ03GiuVvk4db8h2q2PEKdcoeFT0o6AJQX4MS+Y9JLT+59k
sQcYMHzrzCEao0ug4X/YDby54PpUKAL7+CNrPfiA6sU6g/FFBKSdDDzKYQGxVhG/dklpKUY7oC6r
vhr+0Sk/vq+2N5vDf0wwpdxwwGPhkRWySiPx2kV4ZNEFNjPADy5DZ9lkTfRvHvdMPo3mXDq2XopA
R2d5FuLPU1wigmm3jbFEyl493ROVTpZdMncvUZDj3UQBpKHzxpB7H+oeavqpjhKqYNkU02gmlRuF
2xqniJTHtVXxJw6YsD86tVkb1l9rJKVNyzK87YAe+05iy4aToo41Un6Ii4a9W+L/CmX3mPwIBuwz
+pZdeh3qp5NTyzSYu+qUylX6Qo3CMA5DheS01EuMrhFYF/C2KjAtrP9wqFFZ/FiXdKoX09Qof6tO
kWlvrAT2ZkSjnwVZtaGmavDVa2/xYfiIUdpt/uPD/Sls6eSHGVWbDEXdDYitV3aYzyBHOpoWKn3d
OkD1S6q/To91Ykwjv5nOShNHvRDP32jGhggP5RQb3RijhpjH7NLGcaSPtPPoX+UQ+hCzjU+u44iE
n7f2b8site5B8cxneVcwTmJUItCzykpLmOmeJSJ/A/8FnROU58AAR/B2i5mk6pMTrHGb43J+SS1O
EqIUQtIxx7EjCy3XUl1GPYOswmV/ZV2nPQsueOVsWl8hAQyNq7QGeXlDil0zydOanK3t9DTYcPgI
P6iSOYBB1MaVVX0mtX4DBPUnTCenDhts0EHdNkIiTVUYI/2/C5RklBzBQyznggKSPwyczPlqpfO5
RhHVeeVA669m8fQRaEdp6oEUSIM3CdiVF1RLifjd7Ua0fCjGGQfi1s0lvIOjY5lHZY1oBmOegHxZ
gOVc1m+hOtipDwOZXOYe6x6YmgV9Pbpk3cjY627RyTGeMM9EBI/ptJwHYVZ2/Fn2nHRAgKNbjXMx
2iRAE/kc4HNBT6FaLsSFbkji85L0USDDck6l3+xikQLbZfK2Hew1RpU4dDsI6Dwimf1YrRcnliVg
xUGcAYkQDF8uiXxcwowONO8zcfItGUl18fFWlhp2QuTVepQjIKZcqqbeKYGTXFehGLsuhK8vO3rw
nEux5BtNAFtEsA1gBI8Hm6J5Svztq9Tu9voOwV4auKHATpPK4XD/ZMxhK1Y6Lz9Ew1o8unQT1eLS
Rjmpgb1qzQ8KIn2sXFMmRZ+NoVQT+W5ganFMGBMQIqg3g/7ixmcmWEuhKXwunzFNUIUsrnzpcx4T
LtjNiN8ySZbdkVj9QpFNzptIkcDk5sSBnKlOiYZf2RjHc0F5T5hZaYhfA4ftdA6qseLwWftqeX8x
vW9mhHIuIrZCDo0uQD7Hj9Qb4Y43porU2DfHBqLGnb4pP1WSTMsiS/B7awQdAwsZDUMXn4lEJ9dT
U++aAzYNI/c6zgwwAFnUM5p2v8xTBvow7v/8NT0fSzvthOl2FMLyOLDTD5pK9IoH+fhB7EZDGK8m
V2krxIsXcIcFV+oOKe5zGR5SV2en78D8WSUSEf2XrWuq02GdgZuAIQ3GcqSJHAuUDDaefxGN9UBZ
vgxBMZABX/IEOqpkZt16AMu8RJat2VbhxejN1Bue2HWZ69wme0dmJmRfOzthmGUfMTzNsIdSAiL4
ZwUfTmJftzpCJv3FqRQ3FOb3rWVGchhkvYCpGIKyQkai5liVMac18zIjWdU5uGg3olT+67EEchHb
c3QqcQk1HO/5hOQBYgPHUBas+ZZYwq1M/6r40GC9k/UCiN8jf7Ni+/oyGdb+0L0QbnoY3ovFN+fO
3pZyWOsPTrJvnFw0+mhoBa1DYhHSZmcHDegskDqlrMKyQ2pGViZ0nkIKOunQlZ69EqdxnKRIqcOF
PuNtexU0KzGOrKVn6QQipDoGjQh0oN3Db7EXR8ZsYk4q/Zu1+o52nE8jq+LJD5dOEPWdRCN0reG2
pSFeLow+NPpBd9Bf2yeFfDvqQGAy1mNarvrTdmYpst6SBP4ZgXNEtA+qV3iMnzEEDjDY//646YqO
JUskISe+ckjkBh8HvU94eabGKY9PKqOXr6qjoxE61Me7ddvb/f5uTK6f5TeNgqkTv4stKlvQIsmB
4qM4eWtRCMdsS+tlAyl8fQpqtiwnScrY6GJKnLqEiGnBZIaFgxobvXCzZia3WSRFQDekBcRkoC0N
TW6pNRx1woUGKLRrUwQm0X7bhvATH8OPuCMJ+X07NKFfPfC84EOaieaX9U9yiUZhM80FRzV+DPKa
yhzgjrbeHNPaL52Yh0Fe6BgNE+jdJA0+QDNF0tbvAarAsZWEwdWG+T1U9niCAF9hoE5h8SAL+987
IIjelM+3H2xnkski0sg93HHPKDZAu0hkzW7ekX9ayckjJP76x59queOh8ZrAy/0BzjwUOKgUdVBs
tmWMpM6y2zErvXkVUMsqP7Y6Y5ziZMmJXnsLrlyRKIXLYGEp3jy9qBV61uhp49p7NwuKVy4F0eeA
Ne03KtbPs6AoUI4jouEVTbaI6u5ek3sbbKjYOjgUm6LeR3SYawqsI04iVn1zvzFp2wG77SE79CFS
PKcOwkwLIfi9ng7lAETqqz5Xfmc6x93ozrxLhOS7e60GOaTHPmHmEs3beYu1lGr7Q0/aHR5y7CAM
0Vl14SqDbKAbPmjbmLAPC31ygJtNjJgVke1ze8IkjTjcBE2fe5sCUsDCIZiR/U/7cgMVKA8ulDLw
/UVZW0DuY/q4Qtp1fj4TxIt7lOYMcdzVwwrn0TMots+SSbA7l7W/DkAIfWQwfKF4h2rWMihjW3DX
AJFDbC/Wu998mNlTjIXf93KjiRlEPbxfL5H7qAluoYGlowqZaK92ayiftnojSdq5a5al7mUAtv75
YHtxpnARBIUWLM5thcEMBsBlfG8zEYtTgvW/gcO8DjcV3bPvp0S8kQ/ncSdbG3MMgq46szKV3c4J
72LXpwB++O4Yd7nZ9y4unn5cPPJ/s8e6SFPnBaU9opTkOvGdW7KHALZ2fb2ZjzKvg2iZLR+U/U8Q
2CMrQO+LHfzUkxnUT7MNSQIeZ6N2Ym2WsyVTYHY86E8nog5mTzKrZ8nz4H+kGYw+RjLlCtYgMVDH
ic7LWJ3yvNXuGxm7tI4NF0fu4yueHPWH7Z3y7eQiU57ohscCx3+M3S92gjCwA3XECO0a0jnt3Gnk
DIv5LE2aMeRTKurUCz0zHjYReTCfra3pNqhfsyJ5lYGx7P2VH2As0INM/dpwqhbm/PRTfU4wvOE9
nw7aBifAZQyBU2FAyBfsTjvEDwTSdssVfHt/tVW9jrjH3c66jxdS6QJ6KYf2yqU8IHVhKJ6cBjX0
Mdwv0kJqcLXHKSiNVdPC86SnzPBWxgnB9yAnQEo44MYiTZHTcWbX8v4+XcjC3tcuvqzSEF8hL+e3
Ic0DefKVFyWDAZ77q3YragKT0b2Frb5oJKD+vmpHzUsCdesOQf21z6kyPVs4QTPp8p82R0P0Ji1a
DS0wWxS//VGtOd2Vyglx7ly1Lx1XXjxS35j7tyFLBUQdNUD1n/znuiWwnsq0OMKsZR1xvhrnCnCL
GQVVRJwm+lJtoS8BebCJv0lppnXqM5WD1f+vDnSHJGMydSMfeV1HYN1ScMpQfN63bzqrzNdqWkPs
jL1PRN9mk1N1oKhXxN/8v9FCwbjdUdmjBX6CTScrn4uisU+wsfi3l3icJX4/ET2QZKWLRTxLFg+V
nRoSMXGnDjs0BCAm4l3qIhxisk4pKw7/LBmdDvlqed6B5BtyeIGYc+9S4nAsYSQM3KOZAndGj/lS
jJ7SqZyaAGtOo0PHiS9p6I6ov+beK6LWUkwRamwNMefNTwNon7CntWkUC0/+F/8JWDIHVDqfkMO/
8Z8RkuR2OuetcG1J71pQaSxQxMcWLHwNLtHG0xXPFwfO7XseElv4W6WunqemMASawDS0TsG9CUcY
HezKPZcp+WHL0JPjTUgln2VGE0kpV67xA/Hn42k6B2YuW/YO1UqmG23eqR76wEBNBEA5hJRxfUrZ
NA+0FBRiPqB70e3+k9rUaQsw1c4h5lGqjE9U8ct/coALXoIS6aTpVpmd2MW+P1M4KTOrlbGc7KEr
0RDqHxvYhjDwLdHvKZd9H0rz0ger3T4vI1idXq3HTwxZcy91YjSmxBM9BNlvkvN13P8rSIrkPIDh
2FJ2P5Imd2tvo9hQVMmu3tSxa4FBT51ticDV3c6VP06ygAXOfYuI1ISM/2P5tmjFnugF9ScE/sr0
HJ1EQIFV+eukrw9IxADqEPp1y9w3lXWSHiq6LQliUXyN2ZzQits7CVnnwA6KKK9ce9G1nRue+n4N
WGUqJTmPf0CBBo5k9fMl1AdEiolFoCyIAU1rGccwsKp2vU5LzdCvk2RfLJj/fgdRGN1aIRBR2TUg
ZFI+sbtRYUN6igF9q3LTiHaDINlRq7koRZuHZ0Ug1z/CAOupwsc3rad207KztoT2Es3EYZeG5pbq
Cz2N3iJ04yxllNeFUi8HyfUN9KmxdrfT8sA23tjJDatRLzBRE56w+BMkd6YiNSUhK0zZ5RM9nGSW
BN1WLv9CHHD1GnerJyWG0Pds0skjy8VVzwnygdMkhHMnfMfD1DP+6a9JW1pQm71Q+B8Ar6ZKp7YP
rGW6Ey7j/MabKNT0Km0gln4i4l4riLaGjaiDN9jmQ3uvsgnvYZErEIS7KBn3pQihNqwAdlhWntdy
6oZxJkjacbqS0/+lmfAtbznC3e2fDnestntLWIepTuajFYUZtdpehck+WhQGJLbBanCZ1PmQWumG
T69oAFLnrGcSWPlSPl6ozspZZXx/2opOJTLetSNfjhTZ4EZz4AVliiiZOx1SDrfYGvX6E+u1Smer
H2tX+10YJmdsE78nq82odX44pb39WwakV/Wo0bsUtyPe+WUpsmagkiP/WPjlJeyA7ykjZaWKW64/
m+42onzky4S8oCaXA+nYOsEUKEamu0YTq42yPGod+V6LYv/VIhennQqxqYGJdP9mDgSTTiaFBfeA
mazLyBugSMLN+801zVUsZHinNnHPAKZXQsXVb+FF/+I3daloX8QsHcQSgRCr7Ip4ucl/9dyXWprT
IBamFyhDZghHi9cYuaq94LiHbAk6wfl30uyy7F25aaIm9QnHwLYhMiqjDzbDHUTQQBH5jtduVf/G
zrcm15fecbjQSOueuhN7JNmYTHe7zS54BrGeZj0P1Iw/qWjrl2HE/bATAJZ6hxcGS0XUpU29Y3H6
W7EJvSXWozbAwboB7x9xAmQ1sUTADbxR4zB+L+VK1akWt3AE+peW5pESiEMUFmxqKXB9QOHWhxBF
zq3cEv6K3sDrFSeWok6tULhpFhEf+3Xxlva8WXYjbEGurtmFizp49cqUfGFRWyfHOcU+WeJL6DnS
/NSFe/i92HfRrUksRRxDClxgoj+Iy0oFp2qcJ3IMM8/QBDuZGNlIxMFizfzu8c0R10XI3SfuDekJ
UejFnl4jXmDIA/Exu72r+oD26s2UdUB0v6mwLEUV08K6Eq4Nxic2cet4pZarPQVDP42MZ34byZVS
kEyiEIvjNBb0d3qIyW8uFMTCiv954wGMbhnsGeXz3EpdTnqcQbKucTxT1S1pJX/PUXiRXe4YiKdC
TuRgrC9O/5b9+mD8U9+B4/wP5ac/pjLs2EkPPmrNWMsLns3t6rTU4tS6A9GWSShltCduixz5p5vL
/GKi6KZSJWU1gcV3jI+YK3CGhjyncB8o3fw4+rylyD2cOxg/x/Z51T3iTUvZrGE/Fsye+2Ju+t2d
8mk7dH+S9KhWdQDN49O5yBqEYNtWUOeCwXtg3/yhJrR6KhcIWVddmtJXSsrSiznxww2a0f6KXRdh
MscsQRhPZfWuYjkIGLELcucQb9ffquUdbyRDCLUhyzpB7U5A2Tt24WkI4LKfv/+lpr3B4LezDRQP
XfHjbkTY8wsaJm0ru9POS9c/ZryjX4sDfDg/awaG8rym4Y/9IaA+lBM6UU5dnNp/5gQTptEW8mNN
b+drD6i1HfQKv667kNKoVPf383IXuAPCznU1vwQa7a05gX7TFqbLGu3YH131XUxTKtVabiOUEzcZ
RYhpHsd4seSzTFL5P4MeXZkpvlB9XkkJJsPhOowW/vn1bCnKlC+RDAeY+YtAvbM+OdDU2xcnHZUc
7XAWJZNENA8Urjb2av5Fct5Np6j807dvlHNSxo88Ug+/3x2K8NyAOU4piNv4EcpAZB5R5/ZnpM6J
9wWo0rAqNK3tiwnZ1XlgXsxiuc+zivLeH1MrpNzT5DD+BUY+Y3LONWc2V80IEWw4yeSDvl2WNSrk
uptE4h2ZpI/Q5FnaRvOI/JygmamRipfEw5RhMo3ldMyuu/ioWfbNl1Gag40qoV/I00QI4TCnu7J9
oSsDyOcDuyQn3ubtkrJ/UjKnd98EQqBrSu23n+ZFVJEfAduHBVmMuY+fGkdIalfjLmlrCBtVEzp/
PTa6Isugd6qhXEnK/lygLUPiXDV2VJ+oYfnC7bDIZMTHeQv76a9yRmpgNRjUWxZ9TxPlQaQDQ0Ow
NnXXnp/+fuvNB/GPEbHB7DpZmQmrY9S4qSOU2s2oQOuQmcSjLag4Y9ctCtrHxAJHLRE0hb+aorPJ
mgLZO0oS51np3ti87gkqVRt7HbHByynVXCrD7++lLLttAOQzEo9jzvjJtOrgvMc+Fsy6/8Dplz4m
NieO56PCrARO7QBsIuq0ec1tFjVnTmuexz9r6getuGTYHSvfdQrD56xD37Ei3QWM+6aFTFNPp5sn
eNlE9x+7fDph/FiOZCdKmfRDbXS0OAtmJtjOlyAMGXJZHQ1sadAecOPrKikJ7VJST7y1KKzVLjx1
5tLu+yaFzgYdYZo/qAB/fWLGBn0A7+UhpM5Lk4E1NDCEWihKn7JgomeKEy/opb6DusJ0GJVboEt/
qnoGX4rj/arsfwU2o3xbDcCmtj0jQsqdzDZ43MzkSKGie0wB6c4o9BcPq0OFJJmM2OzutSSj0B4K
DH06obaSx42YER2q0vMfxnx+SYYJKrdiXH1KWepjQnkWq6e1yhhyoZRu8YzXRv+HiSiA79YRqLQA
Yr1hFWSyJD/Q7gtcpnd3DOg15k24F+mAZbv+/M4dDDd4tSCA2AluILFAU3y/kJiN5xiAv0fO8Vuy
KoBe3M7/rJqgK4aNfzHXGFrjHQu5PuMpOhE8nYLDdqoiQY4F3DyLF6u1eW9+/njtjN40bM+WsuQ4
WDOkpXE4HyyysjqFd6xMenBV2l7Y5MvHKt6t7zuueWHTDnqpva6Ji+5NgckcL7lSbfliUY/HoIbq
B4TxjXlrsC4sOxXQ2NXigrVMXYR3XyiJCePRth3E2HQ1xCkr7SHvGAqI+JAZSl6kCJ8OhdM7+8Gh
RDUWFI/X5QQy5gL0lJMfMk0JRDiJqBG9vBekMIZYgz1+1LJmd7C0kyMWFu9ts3i+BrCpDQajdLsb
UDb/sXwibcoGUQzOVPMMOpvQ+xEfxirjX6nw5ZF1NfwnxFHNAFGjUCIIFBBwuYaA0HZItokGtuY9
9RL84yPpThCTDrM13/4COl+MB4qyAFP1IPJ9jB/oQCwBSktnzxJDSGU3f5MoTeanwsDrvAtVTLKe
QZcjD4+9Fq63UovfXKORjfOp69ydEVHostwYc0KXHx+PrWSGFYZdRmoh30ENi/JyJRSpTsa8/RtE
uGv5UvxwtywGQ/XVIdaPJRdgNGBtt9PIR9JGedzReNFQ/YL1zMZTNc3uYeVvM0uSJj7yeUyTTJJz
wbHv4Oyz0z951+9IdHgMvG78qDD0+wyQb4zYZLlUaTVp4xNit/mRlul0rxcL4tftKXU/ypKZ0tPu
gUp9Lf0VPRDPVy2ZX8H5s7R0G4U7v3usfKviPHwOOPyMbGG30RlrxMWNyiTGdQJqFe6+i8Ll/1W1
ydLVL0YY67ttHBlQvW9qe3jmTgLJ/bkLmF2MiUyVbC00b8KEbs2FAFcPtc/wEu5nx42ztd2OI+xo
JD74Uh3yS02y4zkV5pnoOy4wmkyY9Ii5s41dxrljBBzp1NQ9ZylV+j9BfqRu5+V7gtaXq7PEeG3S
hBzk+wjpkPGY+LR8Plj+HcSPwggUobP/np8xAZgjFZekgB5pAVZZ33apvnBWW48bn6aB/atKTcIz
+fxO/7CVujvQn6Q8K5NNOekhEq2jUgHfzIMmFzNHofArvfK2VzxeAYrFtj5m5Fa7QVhjMlWAniZV
Zz6WhPpbcvM2pobHOhJSI1CPAbxceI2Kf/F9FhmdDe0usjpiPkOlv/SY/RAhmebMvzH4ODD8YAWN
xrrznJ7rrJylAb1/XuUZtRs+9u5Og2kZn9+t9U64v5GVDOTlFfzEvGvmWz8X6A7ZbjcYzg6JDAbx
fOaRltZ4cdpuvz2VVv5R6rnGJNujKNFX23DzSWCaps7ECBh9Mjk27uDeIK7aCRlJmERkRxx0++tF
VPTb4Tz2p1XLhH8WYeSkpjA2O6o/jXHGokVlcr4dwAw2R/QAc93/RvT+mgKACn9XPYNLMddC1izp
HPVdcOfjudrCBLR8EO6unJa1nNpKBL9R0rcesHCZTaoAMGmPTXF/X4sxMmCenCSw3BN7IhaXs+md
Gz6sNC8HSI8ccp7lhlKmxd2thbWUXjWyQmOd1WmesQ+Pq5HnFoj/MXZ4RUN0jTtrAOLER50ww1u0
fQESrPSgLH2bf5xVas+9v1Bk0PQlIDHBQFn4VbuCBlepNWOrK4EpVV5TI2hCCA986HZGi3xb/Crq
HhrRylx2kT2WWLGgXTOR9qOxJZEVvmL93xCkMn9tiNrUMAUO9DaqLxwkT0Tf89x+uuixp+87t7r2
41LbN55QnAQxqonm5aUH+0XBbF6QmRn7eGx6ay/awdbF2t1wRccM4zA/pL5VloYg3BSclU5Ss0iy
kBcZsxg1eOC9QS9JGGgCNWLM8HJiIT7GImnDV5NNnaker4l2KpCNieFqq9khCelmMiN1Nccc9FBW
CAFvAvCtRIfwfLhEmY1FESGnFby+cGLQomv0xNjxFRlWc1ijOgFMMPoMyGwAlMUquKvBz6svMCIq
/6mTcrKbbdvqy4arOEQz0apy0OWBGzQYMKGejLHoZrPQCJPbTJMqJqHtXQzuvKAH3HoUoK3ue+71
JJ8nRd7iaxIWsXPj18NBH2QIgebHdS6d0nX1r1itIEThuKGlmoD2DNyqCGQ+Bem6KjmU+dw3QLEv
3sjVDeSGOdcwMJAGx+TwoMP3IUl1HYIxH9V7q24RR8LMOK/psnOuPDkvoaznAQJEB6Ayf+HjOPk1
kagPkMefV2Ns3Ex5mRRW3xbJJIY7kJLK00B9RYVtjhe1a5PDhxrdZuNzfI8SWekr02Zgjou03HKP
TyqfFVMZMaC+U6YkWjnvOS/m0zqN3FZKnczzXNsb9eP9CSbZ3RXCIy+xgzDo/A89wuo0yZ6lG3Nl
38hzZpsL6wcRu+8L2CLRuYjhyHVVZJ3a0n8NzAaJVYzIkLFV5CGIscC6OqOuO+DH/wITCag0HPrZ
8l1qOPgR0Ziaqqu3IqTe0hCPWie5y7+WiVPfWWPuTHB2PPVIQABUnfWayezhpsLoW9CyoGgoSaug
Bp6SHEHvqUSbcmhNZaZwi3yBN1OPBCUrjhPNEA4jUAvwxItsRmVMQMegiqAZwfLfD8PFLS/y5KY1
TnNtSTWcWyHyoiFzHC7r6dp398jmO2bdaQm30rvr4SvTJykiJpF3MsX8VoInkqBG21zQAzDDrQOp
CGrg327P2ZFcbZJ8xy2a8P9cLeNjZcDtm4G/eCn087PfrPgfN7+PGsc0PglEGMZcu4Tkr2pbjtfE
5uH8OWvSzZBaa5EDBsk3krYLt9xDlYdjvpF0ptprGdjFx4nC0htC8WhUt4zZeW8BgIabHIjn3jJX
rwsgMDvvT65UfvwcwkBRumwzFV0EFt8owO5zwSvssridjVufY+jL9fi4sFKqG0vqxY6HLyCaMnr+
1aZ7hLWGi61ObGcQ/NAp0LhBy/bFCxbAlP9EJviaH4S1RerCC4mSCkO5mxvq/xZyGV/waIq3ZfS0
FTW1nkVa+WeT+WFj3vbu0NCSUnCmT6pSaIL+/coI2yFG0KX5uZbF8pxFV47TmBF/Gs5eMVYzG847
D/P/agEr6figfb+HcAWj62zutrXmS94IxoeoCGJVfnhluH1aqLi6OrmryJOEu85x0YY45G619UtS
lZfyukIW1BsEsPOZmPqT9aei4w4sxe06f4ivYOF8NIL4GOhV9GHJEBexoCn1G2zpiDPbk9DAqJeX
+s+HVGZlemKgYa0HtlbRjayo+/p10p0NmyvbcNzH1InKiSFHA3Ifvngb8vUIfr0YR/Wh1Z+/QADF
DYunztbOUAx/nlALs7TBlaTC0bHdANkgNCaDuXwuKrEsnRFiBs7aDyQi3OIT0/jcrlHpWpJINVPv
9iokkc/ZcE9UussjPfZAiKHDXUqzobpmehl1U0mgb2jznMKLgmuZ7igYnuEVAAj1nXS//QuD+VCj
OFPUtyiwere9wCec6b1C3a87h440ZuNmz76e+0p2nDujeu2/B1vS8tdv8o4ZAeRKdBi/4hb5P4zM
PEy11NxnDUPvucnHp7LYI7hYKRj52EoUeYrvrzT0TIEWUuWb4FReSKVkQkVUv4OPYEuw1SlrdADD
Hdokkp7Z33TdmtWYOJNIQnNxBDoPg+DTWaIblDvQOYXmqB7XViM1FxyTmNw4YgtQoVYFvYpM689E
2NIbUvcVN2JYizZhK0wAq/mzNpMC6hZV2EpMC/p3SpKJ7+Otgcd//NYJgfUCU6M53mq0QcMyrpj9
lN5ogQulTdRRkI7dbO1KADiiNjSN0XJgv8Q1GrJda98wjdm/Mu0QT/rNu1JGEsyZM5R65R66iWqv
551DtvqVa9fkakngnGDxFI1YgbBA7JNOQFOGXqQk/BcWG9YlzCIqklcjKlJp3OUVyPvyxblXXc+R
3wF8F6RkL/W859ULnE9wvCtC7SNvpQrZdh9kDnFUiUoK1VeF58V3dMHx6VxxDMarTx6rgNKnFQ3F
I7Z96koFq7DQXnKRyb1UJZTsVyzhp/gsrW4inqQQilyJGxXtahuS8ah0dPeEItZSOOK8gnVnLdki
qCknR+r4a32pxQpla8m/nRPSd91/drdZdpOh31RWHIoGvn0G891KNuTyppKxHAjvOU6+biHrOesV
AdIUQkpss/sSX3qkH7lcQzWL3adNoLo+t6WuoLhL7hZzDQr9cUcP05zZHhsCeFpujxsf+KTAbmyh
9hLOQQwXp3TM4Gye5sJGNYnwFZW1oIevl758KB8b/BLROQHuuxLvDtqN3+7jJ+UCCaqvYfAEx7Fi
V3aCjpG6GQ8M0p3crNbGrPROhsZyEgoIizeKd7yudZ9ejp7FnaWp43KZg5iRpDW8+ZWLuVysnsQl
7Gxcml1OfDmwoe30m0T7+f4zMv8ZD8qeshiJQB1gTfNcT3uM1Wt0BVY7NNgFhfjMooBJadFalFsF
b5P7jZuDf/thOvWnISU2Sxu9B1cgNmBJTMi6eCxuiB0c+Gq7aJeK9rFE5r1DZ5puoxuAn5uI1OrP
7buIwSufW8Wk4fWt0cpLQMFurVMAiLL2aKZ5lJJeKMv1Habn21Z5lIBb2gUy9i2oQVIHanQpHQoG
uibuj4f+8dOrQ8Mi58yXxWwNcBCW5+WBzh/UjfNnoiQASnebu3q84g58lq93uHKBGJECxeE5GQ7t
m2f+2H6QPAiptffr+pzZ5dy4uIWqe7ThMC0TfCmf0I/0hFvVsUvgh0hB4j4vdMP9D/TbwKVDzAzB
PsvHWIq/z4642YiFLtjZylq+Ij+ZhOrjQ8s/FMoTmqDF9MlN4gA5paAoFLlYt1mXqRiXXGnsCNuh
AJWa2lKmfv0Hhz1g8BaKoRrt+2uBLdxoH1PRncKiHC4HpG6lw4Zz7kmerrMKZ4x2W56CzeOj17d1
aYOCfP6r1dSG/OXYBuNQaNm/KugbOpUizjeEjv79cDTn6KiNwqAkPy8ThnaeR6B2aEAQTbq7t5F5
zF9BcT5u+/wJi/diQP83q+VajI2LwJRpzdkzoWMIHskL9C3q4ZJFcYAnFgS0rncOoUeMnwnpF4kU
MebEqmMVd+Wjmode/CqCVOMLRwBHruhjgB6488bucXPAWA0rPcMpKdc50QZ0KUOviiDcK9752B5X
KCO3wM4Rae+GmYmo/v+kxfeCNV2WPhgPzA3IVTp7hCi8SbT+AJHhsKZItk0es/tSK88vtPBh4bCT
vSODM4nQ9zFqh0+nCj6b6qXIfKK2ZEDLio5zggBs9OiCvcSD+e0dKLsYNmTVxhaunYod6sBqX93o
kvaHKD8zr2s8QFAOkuKK+kIwAseowwExZ8W4eXRolEYpsF4/mNk/s5r6VyAfuCpSloFq1hA9wZ71
hkLQ6BJL7qRiixwwMKHWshfpSB/wNXi5eVsWuRwFFd6q63vaU44kSKhFmwbvCWuTIRpa38KJQ0Rj
1uaKObqkxuKOABEjuRDRWngNOzCKcWgS3Qo4lPy3AvVCKjQQqQmPzWkBcDKupiIogoDOP1RfGmO/
+PyRPnuGwZD79ixeg7s78yFEnyxuMGPvG4LOd0aAv70hUKhchXoANxsL8UgkZcD1KQ8/rmrSJLzU
M6WzMfrx1cYx4pPIUpcBtWE7fAVqwh27D/XMVijV1ZzzLbgjds+JjFmrVpxUDPYuxX8C5ShrOJDc
DYxNh/IRWZnoMnGNuNmZQMLpDXrmbnt7URpk4/33bdacNRtt+8iYimuZDUkuGx8p7k2vLGmGK4mU
gsCr0Dwldzur0dJDuVpmCr+S136mRz4gWxkj6czJ/R11Ze9GuAzVdqhgIU4xrZlH4Jy1ZViQu1MA
J3gF+/AnbvmkbvgOc3q/JdE/VTqiMn7KW2OJLpC31v7LbZbo3RrN30TaXAe1yr4LnwAANldiIO+r
wj2h5+nJITQHELr7iwu2KGLArNzZw3A4BTUXqT09Rq+9S+d4hyrYYGsVgResrLzoqOaURs3ReQW4
maTo8wR086c74GgJiF1Z4BzXTGvfPJxhw9KCz23K2u9AkUOq9jh9OEfNjMLLC0Kpua6Vzm/m4sd9
yVJX64VjWNOFMPkhkM5TfqaGr2Mz9Zv0Pww91L3Mebgg+YA5FAL7p+BpJooTXcMXE4wk1mnQk9YF
zxJCVGGl21TGkekN1TqBGoku2srIsg5uSTBObz9KehH+Xnz335QHnGBlE/hposcAQL/snawNBjwJ
lCOVqN/vjJJ7yLhJ2Zrn4qAe0pV3TzukUpVRhPVK+lXNoejo3Uk35s3dAKzbj3jXu9ubY+tnmt6P
zmcxAvAkx8AcxtEznmkUzQhAlnSKvA54pRVOEoMGdk+kV4yg9jNHSega8Uhpyh6zawLxhRVs/sUu
D1WKHpn+7DqO0PSzXiGaMF/11B/lB54QWSnz99gzYBE1LAVlly1BhO/3Nan+wVpYuL4fBdM85TwH
doLdvac95r0sr3hAl4tPT5hsgH879ViL1ls1h7WhWlClHcO9JjF/AbTaR6/Ei515aJ2g5YxBJiJL
pOtUQiX5Bnd8qDyGPh7Srrh9wPnIsgik0xa3SZ0KlwA9opYpuKtayzzMx5QzmLWRsD63Z/tm3A5p
+R4DxgIQ3MufHrdz5I4RmqILs96zo/K3a8LCGl4m0+gddzyBf1BySIfj5/SZwOwKL5UAquY89JG9
2HqyjC22e4E66lZyz0hKFPLQGtuVuDwLxxO2VAqAZENdG9e8VV8tLtRMMHJc2+GPCduYUb8/hsT3
9U5yO/wAJFH0TZayTRF+6Qzvi5gz/GwNNljt2miLgsFkNxtd4UGzipJhf8q4pALI+NobTzH5VMTg
jEnHlypK81HTvr3MrJPUV1CeOhZcZWMIUMTqLaRSu+COKiegP5fUpd6LNr0FAnO9ErO/dCBkBEYR
I9NftoJz9RRhT29HRJ8Y2l81w+Xtc4S4xD1efCDHWPNudAlaCYnMsuUvKC6iKUpB8xB/z/KsXeYI
Bl8Ue5/ZCVo8nElWJv70u8vgllj+ZuQLBsoN5VPwaXYeTJA0bAfKhjNwymyF1HoGw5yyDeJl5EXv
+uI8Q+lztpuSlP3gychbvkK5p8KfrYUx6kuGRhljOAPXkq89hXrXEblmPWgti6J9OD/gJSo7ZCdp
2LJPmIa8bYTKHsYKAiOAlszx0vKv/aayWBihU4xQKAQDqjlkO0D/wKAUBcnDi26scmBAjr4v97Yx
jPoOkswK0HFwu6fzFNLAMw8mvkzQDNED7waK22yht06UDg3IP0IGrYP6YPyez6tfreMgz6n4Ha4K
RJ1o/ln585b1znPiGqP/UOiR2UfKfztsq1kcWc5jYiyMy8XV7LLE8E5Igo1AOPmLYJY8lbXaOGry
Ug1aCYdsSfjiQR2xtu9o1tyQcH6YuGO1HJC/qDlqDDP4ngN2vyqAmoncRFH9o2gM51knVtPIhMey
3jmKyNh4xx0odFfftoOBRy6iZ+oaifIq3z5kXimJ1TOggX+l8wuYxKUyEA3IR2dHP/WPM25U7rVC
j0q3oieMwEWWt3+t2kBZaqCsohfj8gwSFa+1IDe/2pHchr5owUf6tY3NsBHONTBZT16fyy9ZURcJ
tjePjJ6IMC9qiN++gwY1ePZVPPBAtF4I2Azc9mjQOHKPZrbtEqnGjubtRlAdzkwf0Ca8M8aejERg
Vdvki9IkG+n1vyec9qOqL89tgqrKkPNOVxV0h/PmaLp5qQtB9ncy5PQ5w5yP04GBmvTYOBz51TnJ
2MA+cH0imqfJm3A80AbPL/nPKR4YpOh0DNgI/xKdwguaSLkUu2wqiJ8P4DWHWa6X3N0q6yAzhO1A
pgYzyZRWr//Q3mqIPFaeqlduotPzxHDQ6ZSd4CemprHxmdCU1EbsEU7d0FIPkTIPLjjBfU+TZC1q
r3/6knjHyHhE5SVcsF8xkyPXZSnr4eIKodIc+GA0QzDlf5w+nsS8u4msYGt6xpQZenZFbvb/5/9j
PhmKpPXCnwJWAuonxz7Qg6MnFGREkvSq2/nDX4P6q/HEQsZTQQPXRZcX9tHulgl49KYsgQzInKen
BA8zFPXmIhusGmF2kWXj3MX7c3yOxD6UOwFWAz/NGvRDLJX29G0MXCLgBFlqOzGyZZr9FffUTmc7
FsN4np3d5P3SnkFkZU1sIBvZPBUKbrxmBL6F5occS4KhTbajRSW+oGJ+ora6EeJPpUaS9Z8Any2b
YX+BseMFWFdCENcJrcoXxlItKJZUNAy58r7hZSewLBYoWCGkkV/CCG7k+RKYoxDZRMjqlFqoK9UU
VnxzQfik7oimVpceZAyh26YB+096vseBNKsgS5c8AouYGOBhgRmzVxw0OQ/g8OM+zEgoQrPzs2EU
05MVBHg3b/pEbk4LVWk/9ped/yTGBganLwSHxhsIjNwkK/+3grHsr3Lh+109FBPQjrfgqw0tqF2+
8GcOS88Yz1pRw1cITyfio3cyyq3+CAckkC6vre+mE+6uaKuqaIGlow6pzi3mSUmJbS92Aw7PSx5T
u7oTzj8Gmz2jZuefqyuPqb29eZa6tODXlpzJqWOGhaa3FEJeW72TymUgXYNXv8yVrl/L50IJJYkf
CFcDBcNLZTwv6e4jJOIX31VeJhJgTrt2Rt+5s6bzwlaKdZATS5qcEkSVdUZGtUx7UGSmQftF+AGL
9nTGvX1UznwcAhP/2895XrqvYkQ+pn/v9pBO+GyGNnghds/KgdyFsKNAGgWFwKgEQpTCnjMeSCe/
uXP+1j5+r1TBP8UMvzWkEkVpdke6VMAldQgpkd40AiGICcrxsj/4mYk05FlvR5L7fKKT9VZ+hshC
GfPvlAD7R15J2snDKijEl63uqoe+Sp9VhzRCwE9Blf5S3SGe9atE1EcDG7j9Of+mL9aS4FqdapUJ
F3y9mtldJ9uMwpuThi3nHZ3VmihOKvDb6g3JCM8KCOHSYwS7GSAnf3TC6MWIk9kTBNEiTK2lSJsW
hPZ3GngtT8EZyAnYELCXEkmYiNVFZqtAyw4yCARMRO8Kd35ZgeIcpBHLehctjMnI7trSHyW08Bt+
7uqvpnozkxFaiGpxaZnsPScgAUJXvZ/5w0Yfi8FOr36ovc7M60BYoetzSO3jBmOW0ObLA56LJHxb
vFkxp65yz9Noo1etIX1BbUmdGX8vP6FeD4Hrd6i89cYKBNFN8ltSLdbDuaBsYo3v6G1ArE2blX+Z
A02WRfQEVjF3U1VODcHAauwO25Tlb6wjY59q4y2rWsszsR3T+YkbqMbdJW6tvSYx6F5aHHjijQgT
K6EqUhklV9ZrrIlA0gaBGOABMwy1wOw8zI4xBjuJTAPpNxX8HFl5Kawl7x9eoGYAVOIKeCgMP/xP
H9KPwzQMA12bSkQRlLVMWZYJSp4eCETVa/N0V1xbf74E6LasQE1f6ZYwMPb/WNXJeZC4rQlbRwJv
XdNKhIuneYdHybTLS9y2hR6gkpMYwz1fFiDCcX2moL7TCEXaIGX5rArP6iaKiGQMOW/EjSVwJhUV
ih8l12p39tIuGGlqTzRbyptGrKpmecGuFm1p1gElPpkZmYgs8oz3IS7JckF1GnZ1zm2QB/SrMxg1
WuXb0zt8uI+b0OhcmQ3vYx6Wfztlr43QMJasd/gkTV22tPqqRi6qB9rsbD4sk9PynFrm3LMG6x3M
YiUvJQGwWtndDu0ymHoF2Rzx3E1G0u6oZ+DX9DCgObkIbD2Vqsq3jmRn2dFqvTHVUz87Ime76Uiz
Lbj4va0I5wLZh/sW13N6i2ET4ttY5dkskDAsUIm40to+yTTvUGtdvUCIqgpBjT8IYa25HiLfpCx3
7NWgjD3/XHYBprrrivGFzHndk85y/U2Rf3k1GzqB9zG1a6XXOwoTYygNB240McwW+6AwjoddiAeN
U8Jn8DE8SGq8JyE1WjmLzm+vExztx8Mkq5BAU6QFDtvRaVpuqSlTkTM9LKbllMD7v44LgQn7f5BX
hjjG6rzMb1Lg2F+22U4pgErmPonwE5MaTsk5aBVMwTIj3tSUXPA3DvxQWBbx09MtVKuM7gJbW6Zf
Xw0RtkyU4YLYHhK0wYE+EDizqAcff338OHdV4KHyIpGpKNyVrc/9nftPpTGSWyLy3T8trXuczVcc
LYgZI2Xu8vdUqJp6qUro+hlAcKFEXBTvvPXYkR3Ukqm0qK7EIXTvV7K+M0FMBv08kpufawrPguUS
ZRICrDfjOeNJKcCPZJRjDshBjVvFE148KHI/r9DAPvRR51xReGn80LZmc11aHVdo2S/lTthzyjSQ
1N1EPmsM0aa2iOpoP69iHAMsl2UpNp5/gtHQosk2HZIPMhszw8JUFuNWCy4EjLX9/ls/+4n2M6X5
BMWlLoQFrEMytFCY67lr4Pg94LtFYl5+rPoJfAd5m0QI2T65buk/0zjDC8scF+PV24S2OvXirYF1
LbChTWPGffN93dcygaze+Mp/Agh9tvM+QqCQqFI8/QBPTcHutvSbAGhUz9Gr8nw+cer23hAuA43u
XU6GkiUwrfLVFmK1oo1ZU8Qc3EaggPxah3c4y8JiZJXUK1QGfCt54ln8CDYoId90Q3m+JuF0ZQ7M
rhJ+2Y1u7X8SK8OFBAKudAauoj98FxnngFhGyzLvVKft1joc1ArGHbOWlIE5aJ6+ml1VtiL13KEc
9LGBGx8YPLq0b/vC+sFgpZ3uDrK5ZkR8br/wItqTKou2POF7fe0GJqwlNIz3WCBolVdtGu3J6YhQ
uYLVjXaVFGnKhqT4WdGbwSr+uReZOg46GpcDCa4iCNPpqhw7pNDbXrrKmAa4/wKXR3WXrjb3e+6q
+I+F4r1r4U+cZ0VkeKc99lpx2DRQLv3cMUazSoiPcj+FLvp6zfPit9uovTld8yVb/U7dEBgUNeeF
nlXn9TLV1vV2HuIQpYB2cwZWHJ7vFcOiKmnrNqk91MuA1hjEDTwQVIUgrVLtUNoalcGkAQk5oztq
1EZl87d3xE8i4x8ofC/9MMwmMf1+4C8NN8vPW6c+raLsXmsF9zGWQ4TWIM2z5JPEmGwkX3bO9TWJ
dz6hp9TDxzf6no6cw0A3YDy2Tz8WEHc5eYlD0vq1uvddadxXvR3zCbwiTvRc4+M+cJ63/NOXjbs7
VZ0euSAIglBhAJo8MgtocD7/hznLsFY9Z/6CHxICK1q85aNvMh2GrjF2Q6cQ8ULjyKgCCZZRSBHL
hPpuR9ol6HY4appPWWqYOMvydlT9SuxkDFfWWIvGxOM2cEGwf3M2wQsSiNMZp2K9bVMTSnwd5vnf
+3p1EAfeaFyg9255q43KM6skAkkl2yJ22pRo4f0a2gEcaEhTZ91WS6TPHKTgYhvLMEyAFxUBTDCo
3chtFUhI8krhD1tr2qF/lrZYMhem9QUOJln9FXqTl2xux8vTXQDIH4MRrHgUiIcxEy7mPPWp2SS4
kTcHff2ipWyMcIwVm7MTtLo89GwGWxXKptSVwXtw08SpQ/aKHcOusoX+IuBxCm/MjZp54DjnmQqD
8T0L//yEkxAnhFUqbuoeVAXtheXRw9XVUkvHwdlushA+NlUnSkKgpwWio5W8LuJ6t7UqeHTmE3en
0WMDvRZcnR6JoBJY/RZ82LsIfMBsnqhijUBI2ewn3NeAt21lqhZY8+HBcyTm34QF5XRiqf1zjbXa
SCK3QhrNfIlrWJn5lh4kesOs3psay2BlySalBKdn30cakv4K6W9V+UGcwBRMs8htcWbjnHQ/MO+7
tFxx2CCfoAEGfpRA5nY7GtzIDVxSzxflko+rQV8IyKb4vElFUFp8zHVHedqfkz5ZiVEzxmIEofMc
3tQ3vlugAopoYYDuTyJx8td4DJQYrlyXimAyN6nzI23HIH0Xn/IpylgDrU0tnnypsHLEOCxrOovC
mwxRyyuWKa1EoHwzQPhtvpwhgyiNDzWEgwGmdMcjKxyrfI+628UWQced2lzx1dn2vAhQuUX0quc8
Fo4flWOwp4rctxwmNfjq2QefAGpAPBkhNtXX+HTjLH99BgyLIdB64mpPoG43FOAw/umjQGQ2V/Fh
guTDIHyx7hLw8xChsNN7/2VS6tyWBO1iD7jUGiv4IB6rAaD73FVSntVfZuW4nc4g0yttLnN65sji
MZ8n0CfYM4kVuCEZGXYr3JjYJNDe6Hnq39/yC0bw+3QOSYbtEcGRb7JFak5jY0wbLXtErrzAQml9
ogXYPt5xl0qLAbuixCzZx5mWeM8gNHcqGkLhUmQom1LwsbhrGqdUzNlR7mvx7lOjnuHm8vb5iU3z
i8uOWgnIdg/Ymii0zvM/lSYWdpcqc/gZVQgu4zCQfWOpJi5sz3cU1/ZF1MaX23OITJ7jbxCYX3PL
zkdWL4UVihS+U4WgY087f9GI/owFH2Lo9Vmc2XCsPfOGrsIGLiZ7aTbe0HLm+PdVOJyl79GZMLHY
CqgVfioM30cdBNO9HlGIlxCK6RBe80XJZ8IyjDOdSDzryhqAGrIhldYG3ohzjO677iTM7x1auXdh
MCac4Mj6rxUhyCxmMwSkjfIt9xyRko6cjgfiC7FRSNULYKoCHRDyq53H8Pn26zqfFF3QkQGQuTnt
Vi5fqeGQNnyOPYzexLGPIymBScmMqrFnWTos5DavEpZYHNlTTyoesrCBfYLyCc8/KaXHEJTzSwz7
8zKRYjbK8B0IIb9u6dtmDy7A9aQZGXJOf39tjMBrO96tBmvJGrDxlc/97up/j9XNcQCmNZvsbLYe
6ehju6owdmHadkW+v/Jj40oBbDxHycdPDvR/c63pn88w7SeLnaqtYuBmrMgD9qIqVBvB4dYV5x9E
Kg8EYGBZkcsO8qdvTOGsoVjuMl8WgGMX8+TaVMcaX4H8E3Cn1w1XRpnr4MF/tyQRPNWKpXiXWpcT
YTR4hkHqcLwH9HoAaTrc1oBXaKQLxPXXugyI1LQS2ylsy9q4gyd94RGdaEI9XAaZfPdaGNVsPpje
kP/miq8emcvg7FDn6stl0ri2TEFgHs1CpwAq4KYResm5hDCXxscWbdA68yfKdOaHKdYaLBuEVWFh
gkNixiR/jg7yEJICgOrRAYVqASz23vnyFqgXURqpwTbPH6ZeFcRwSkm2prk9mOG8pZ841sYZo5w0
8YbhlN06MGn2sfDq1YuEc43yoDCseKRDgSRLS4I+iYwrbvaXL7WGpbRq7xje1eASON6r8c4PHGfd
OUurGK6TD58YH8BMFkNSAzlMjYDrte5eJMKdzm1CaYL1djoAO6FLOcFk8UAlDVqucb7UDuLRbnCF
/BprweTUzkFha7u6S36IeV39IHUJkpgYXQGpwLgS01oKy/SvJh4qvBkf4m1iWQDwwz9vjlj/QKQk
cH6lUtfuXgMIYEBlTUxQC9OD1hUEm7//auFhFonezMxEOCZa4DhRsVX3cIQ8TOl9JZvEhA8KZf6G
43aJ2W/I7hjpnPK8s39CnvZgNuAvlcyzWogMrddn87bKZoY+QZqWmy72Rq+WSQaWob5Lk5nMTp+F
50IkE5ftWHXSX4358fkR+8cHNCzwanSeX4Qs93R3uio0Vcj6ZQ8m3f6taBldTm37SiqbSmMHYFMg
10yuDCsozyTN+XKyFVjaC/lovcCvtC0vY44rtMJMXsoobwpj67jJFolv8qZdfR0mJah7Op1tnd9D
AbYfwuL7wahDAGvyFsRzLdz+ubUasrES2uXbLwW4+x+gdETIUzpSx9virbyKQKOw2xbedRmLaFzP
icnqbNwyQNcZQkwMLQmbJrO9sJYkTzIWRuMbNXaRckdvAEV8O1O7N8NbyiUFC9tt8RWH0iB5pe83
TeCOikWemeVeBPbUw+n/CADkLdf3ixR8xr3UaeMp1x6Z/ejz/u5vKHVmARPdSYK3Y/tWye8TgkT2
lOibNJLoB6S56ixKH5iaV25j1UdqnmbhtUKu0h5CFe8jQZX8EXQUpV501ebyTF9Fix2ZCnwjVnfE
nRMQr6CTVm/uo3Bla0aDyESixlNvCEfcPRlKCf9d2O1RPHNW2CTAXmjI1xxPKgwvRl4iipFoefrR
tfFStPyOfVEnHlwaXxmH5Pm6wZVG3B8qvRfDZF5R1ItdJ34CwexVTqNaBG1TRsuvfFkwWmqx73H1
T1oYrVkn85I5AMsA+admybfC+ePKcUa5CjN5dHPFmV5KElEHYbNB8Y7pufBk61y3dwUE2y1iGm90
UB8/F9/3fhjP+IemJ9l91MNkDB9ae3h12+CV+fQQDb62dMRSbXS7t5SDYHl4ppGvggONLabO/4aA
RA8sX1Px53j/sEJw1kFS8um2l7xRk7WCLUXc8Qa5PMgtumyoBxwrVMzaQrQj+0QhrwofJ5vMgUv6
qv0Z25OR8X2Ryqio5kG1oEgwViHVCFalOg1U86suW08zopF4T/8Ryois3zmTW7BMF0jJlgRBgE8U
XnSnVByGYQZ3onti93Tvw5K7Y3C7MGTWc/Z0QfIM+MyQHZODH9IIqeCIT31O7jsbQ38oF57Xm2A3
3fvyxyMR1KvBi65tWWmACLoe7pNewUgCKMi2Z5bKlSfkAZxAdnM6TlJxcnvJdlY/O/BokUn6tEud
w7luOBOLrpt6GLXqo5N1QB/JiNdP5Z8AZvjHRrEQNTkZc3wmI00ohlH3SKDvM3A1+Lo9Iz7cXA9G
q77zBd6YRXS+RYtVPR1WqgyRuBtplzxs3bgIv2U0hhWOpyxexwF1r2C041W77nfCsp9kXSe4qvR9
j4rDwiSqdSIYPL7uOZIGWGNTMo7Y93IzAh1T9FAsOqK6f4JaA0C1dGDB2QKhWmFDnEmqlvoacIUA
6rROPPTNDryYg5wP6f46ETyRQPa+TOxlHdeULyB5yA1Ua/w/rLZyb+iMamqBOiMEtooScPXXOnoM
ga0/ttf3p/j+iYrHPFdbgLdfuzLU8FwNdwzgQtnreTONUdSIZ2PgJ2v3Lsrpi0MzLf9BCzTCNmFA
2yf2FfGJqnrqiSDgLfgf11Fh+dwCmAwpm7j2dy5eHeChjhQSRKi0Q2epZTQDr8FGt9SAfWSEZQnm
DwRGMKXmmHgR30O1urDaqDXOvEC2gNY0lTzqtwUxk+BG1rVBEq5BtIqdWPSb4EqTMRGRnDQW3jDD
5aBIKA5hIeboyANLn9fErNylMIWGL/TNdBI9lXoyRiu3bGUaHJ2nfU4+0Hn2Q+kb1HDeLf9WZhqj
TXrPz8X1PB340xTxhpiXhuYNi3QtZUStjTXgGUJRIMKL8kZesLNtf7YZhZv+Px5V1J4NhjuiSS+V
/Ij85sC5+8I6X7I+h62jKZDlmZ2a5iJqS5yIbAkLg47WOYaKrJhBrXcyCXfJfSA78Ta4F+66HfgH
8a/jK5gB6m4hvolrtNuiHXMck3B9irxWiXoFz9dZq55mZbdZmgNXXJz0llQ/yLhlQNWvu7ktSq5C
GaHK75TLaCNmkLv8qLS52C19vIjKLsq5aZJRpuFupJyv+UddGvIkEYFcbSVhT6JH8CcdUzs3M8jz
ApBgKASaaw1yDkhKWYAndfMYkHTerYITL6jL/D4Gvil+yxavzn4/qduA+1EinX7LVssJwblEbrXC
A2Meq98yPstJiwNul3lhvWVcftAHrUie2KApu2kc/TCkkgws7WZOtimy04xtGRIuKPbij3Yh41J7
GetPdA9zb7zPRjOOv9OjZ00Ll+B0CLGle0XFsM/Dz24fhr54OgahTX2rbjU4g5WKkcINqNGaFQZW
mqP+Sd/lTG/UUQSGSRsHwE9/k/RkJBbE4qmcfmb79qdLwVYq6lCmO6nuUqajuXTBW7bw4z2hCGnn
I2FjbjXoC4SBT+4C4bq4HRdLv7d5lMExN2whMqyoDsNEgZDmDIc5AfzGPeCP58nw0H7hoIE2E+U+
bge02NvzIVMKr1OmfqVs94Nby6YHyevkfL9ly11M6TqVzPU4rLem5W8BuI2G8gq6qoLr0zSEtbFH
Y9Y4bCd2/7PFlOpblf7E0gexEX1EWFv2h3n5Zy0rPmHuVdiZccejeJZfYz5sCabSRz6tKbPACNwP
WIVOc8MkzWSntGD4YgxlcsrvA2r557JoKiEWI7dZ0Lkraj76SvM40MCGqLBgIGfdxJYFoT8iafHU
G/9WhPjv/OeWSGkcWFNHoNHs6NjG00sUcz2hEG9X0WTSJLlrVYm1+5PzuktoK164tfjBfBID6m56
Ci4iEDDrlvQz+Ny04Uvvige4DpDPHk8BlTM2XsMS3M6nZfwzQtVey2VzZ71hBeD53tQfdsYQxCFg
oBioxOk4Tra2gjT+JgEuFdiZa3UbrNGWJ23541Z8OYdbC8JYMQZEtXoefpqCMyO2Pfmdh4uoyO9P
PClppip+4pYoHM9sIxQl0ZfzTqIHp3/zU8lgU2WLnJLUTH59T6JG+VzKsOHrharjrkTLT+1OvYSE
WqoKwcctB5oyBAD0t6rs+kUjfoQMlCVGw5Y/g5O2tnFj5GqM0zdcrAyiHSK4XEFCjcbVMy3eUSDX
FD0Uiwci6w/ofSwEuEaXnjsGM7Ns62AyFTj/TAVqeX0BKkOg2+5oOrocvw+SDhafK5MS1skqm+oC
9o4vbeap2KC+18iGhuz2o2Sh6TX/xPII3vdsKyxrCD/tOGlPpo8Ztgmbt6zPCxt2ZzvnlcauoQ1W
RKcQoRpY+77PNkNPOG3AEv7Z7Jih07uwAaCW/N8znuYpsdWiBgxQIbj+/1xA3qWCH3Oy1fX5aSTR
7ZuxEYVsUDiKQ9LWuLNYZd6qF82ogDSH9mj/4PfsWv48w/QmIa+iPYk6CIZpKCodl0QKvgVkveUC
yjsTSFnDFpdWBrldWRsFI1RGPB6DgEhwkSDHze5akn0N/rQTQj+cLjDOfW8fgiw3uJ2dKE6D5uEj
gs3UvM2EpB4FyaghxYkcj42PVwzUsORRvmPBTqHPCS89kKn3GoY2su0zIYAZWILUC/W++m9KpHKS
ERt+28zIRXULJ2FW0WXH7l0aWeRyiAnXK9GZ4lJxBkHMtwMZJ9OLiaCCM7esUE4qj9LQvE8QyjWc
ZnzDgPj+mXu/DTM6CXH2+C96Fxzf6uGb8z+GWzcvHQyEFjTZ0/rBfTuHXiBIF3P6CHcjaVSQA6LL
7bN+xZb6DU9o71dUBkjERDSMVBzqDvidMP8pIEBLMT7PH6uUN3y3wMcDWhQNsT127dUEfHNrF4JT
SYN/PWLoGg4pZDE3o6e5odCwbPvJh6rOckwe1xGhuLaxeR5Oi1gctvqVxr37mnjmoRRAGnEo8gn6
vH/oLHF6quA6QlNMRrUVSCmNMG1M192yudxqaTZumlWUmndyHjaaBLQLRV7RzPbztELZf6Jjndzd
I+gallFirefpZTaXFRuLQQ+asuOuF6MRqyDcxIm1PMrkAV2qi+v9TPnYgkK0OmVqA+CoU8L1WZ3V
OqBuYDfJdjs9qQ82WdVHVHyJM0rrkHW4bVVHZ1MU/e2hsyPEiHpFmAHA/nC5+rhkGtzoq4t9oj7s
+ddDIG3rvfMpbFwoUgx+IOyR+UklHlpDHpuFb4nZrYv638gV4MSzCgn2Ke+FuFQcf5DbaQ7wLGlL
7T0SaICyfXDdBosXRfASH79VPwCkj4ZmzgbSQE/4MKriYHfM04GFU+gzVxb+hiRLCPRUNras6Z7P
GOjCDXJSs7qj5ZkhvwDHhT3i7VYj20qyG+pboUAuw48jDUCfBjxgssizmYTvg4xxADEggNzLp/3p
jyJhx0c/4rIctcCmwk40E8dG57w3a0TyApuPZVS6rJplw0C05dUJ9BN2OuhURBRc5hYFGV8qWbim
H9ulSLE1VpIlOaSFx++WDB1HjeA0NUD6ibyLKLL27BFHIhgvuo4w9MdtpFm1GHcyl9aRU/AI/UfJ
l9xnNXQoSr/8EbC4cmHGapINdxT3eQBnakOK6va794KJ/Ox+Rt5CDOPq6ZWqnbrNS+OnJ7VFru53
W4FjTJSrxeNnVICy/vXTba+jqqfQzr4s+OWkTk//VsdPqQqOvRbMO8wnBCUqJCq9uxL0jp5vlQmx
zbawVtmP+UyUSMTfspWfNFKNBLFzbMYE9HCL4Iqwtfw08xwFjK61ORhLo8UNg5j2HrHOdPHpiSN+
8QH1MV+vntZJ76mySR25Ge6T08eEajw6HaekUIsgjXLnHYxybW46AFOADpL2CZReECboE9ayN/qR
69wt64BIIisa8do1zTvS2Pn8bq9lbxinHJN25N7vo5JNp737uuAXaFdJsR793ga6G7iHMYSGdSxk
w0IUWlbBmt85JWplY7Fgoxwg+2jnViZBn+8xN5mMX+tZ8SB6hycTHFsUb7bkHCDXJiwbklaVBk0o
tgDdh6luxKwkYmdk4CYa18IRsDKl9Z3kvAUDjrEelWN6Yoguhl1YOfoi5tFLF4KhxfvORvgXwq8D
G0ZSBq9a4cR6h7YMH+UbxJ8Ves/tpHLHuEFrL6uLimuqeh4r1V2pHWkJzinxe1wA0AsTPmJiiRzu
3Sjl7OIH2kPUK1dG7odpI1tqEw0bhqZDOBfy6klua+u9Dgka0qo0cIqXPLkLsxxRCxE9Ox0RDFit
W4SNFUOZb4FQYznMTnZRAXT+BE5TaasS+/qheov3fLz1fmFON+xDYtzW1g3N1bPy/23iuHnfEL/4
EIlX/yY95OnOPtTVhoMbOq3eRqRi6kFD+QcZ/aSaRxD6EuZVLd8wW3FD1RP+cHctkz9FAiag1GWQ
JpxYIZc2FLkWZGY5v99+Ysx+RfRZkamO8FILTW7jAYm3hz1ZwG93KmJ4COe8k1OOGsJ2jp6lgVuO
Y9/cVMa4MuyD8xGliVdbUjghdHVdAHbUnOe2ZLFRUPHk647gwag51PA5MA8A1K6vK9HHhBUFCB+l
hrG2YNq9RaJtyRt1WNqhARcaQB84bw7r/gr/n2QDyIG6XURsfrtnQ+qMixpw6j2hrj4Tsyp4uFXv
vjgG87jLnuAw6HWRrKTJKP0mOmst6jV7AAXTk1jBMEFk2HRm+g8BkQD7nlmChsNvffkTaZpLtq7L
ZllWDt4IjvbLOPSpKIQ/HBwn/Fq8Rjnl93qlsqt9hM+fEYjUng9D5hWE46lkeGeqT0iJpO6YL82I
7LlI9P0o6sAT7ZtHQiA+/vXfvzn/T8sQjXmnzkDauHNUVLNco0p/wxW2xQdqs43nVWXi9zR+2nHs
TANUls8pQALeJU+EH0rIomQPrja5CHsYXzuL07+BlqkaKGWEhw4CBYbixtQ1ywDkzlo3mmLkE/j3
KC1KQNkvK8ep7f6KI2NUxCSmHG3mEHj0C05F77y7d/Nfk9FdLhBpxGRX8T0I04q1HFp8GyMAAw7d
g3Wm3J253lJWrdR8rv3hmGpyQf/eETyxaKTcF+ZWtwxUOGDiaj3JwPBjbkrXN5WlfLsnJodwuYP0
ZBiMUaV5GvZKKtOtHE9d9JCvNuEr6x/UEu0NEzUKvQhKMeazO+Lerf2I2c9z0qWnRbO3oaDEctof
BsSxOhK1ILVffA1TDISm3DtXadd02zMaH7hphY+DmhfpLvDta1uIakF5a/7q99hLkX4E8IHweOOw
fePawgwrpJLY7jKeV23JzYFxOd9GZwOYwCyC+ki5QPgu5mkvjRa+T05mVIG0iBx8gSSMR+JrPvY+
VSaiKu+tJzE3wy1rIP6HUUxUdItwspRytV5T6JN95ME/ucbOvN2pOHeRBmL8ZMjyhFmygOYEg7IM
uiLLgzl2VXHPw4FaVLvZvcVttE4m6tZ9DIkMMFlEyh6jTpSOs19v529g/CiPbw2BKkNzVWFNl2N+
pK9tGjjXcGsvCDpvlZgTzHBGh4/81ay0bV/2QK+gUvQdVI+n3r4nN5fA7YYYE3hmFUiIQxPhrLY/
W5jqs4kkuUP35oG56uuDxnTnZAWvs2gnaKHGviZ9C61ayueOL2e6iEj4XYC+6NMtKf4WAsTOiubQ
H8owyIoWxAEctcX7EcaExHUi8LNe+APJ562zoGKfKhM4CfIh0Uf3KQDVXeOfYJcvnlQt2j4L7F4P
DuZdj/DEd5yq4Ysv5+Yy4HJ0BsknDNFvwWOJMsQnMxV4bYA8M9KasgixEIgrFnh1kji3XNV5ri2O
yytufjOo3QnQ6jjVtUZrIcqRfvFOjU4FDM26QfjbEbvUXv3tiD6kccdq9wfHEhOxSyXrJz+NLC+2
GYUvy2cou8HE7cZBb1dVjs/s1+Pg6VVJY35BfAkoZgpzLgcs4swHnqvG+KBZWy2DIyl5iUQRynFI
yPI8el2SniJiOk01gJxjpZyjnAnf2bDIHlh+Ai9i0w0biPjM+0DcNuFc5DzqbVAMir99/L7a4ybr
aTRR2iW7xaj+tlaV5ZVRfPx5OihHCA/x9CSvhFY+QN1irfdD2C1UUr5H85xQ69i+mkDQpTp1q9f/
HlYcMB2U5NrqCnLMhYUBB0EMTz/8FvRWj6mvV01nP3oJkIfb+7zhlv0nMB1ZreQWy20pOhlk2Ebl
c60n4X/Ha+OQJxXko1rXNTCrGmj4dBba7MYuEduwxDwsgBKDj7EWwD76QjmJdJqGlR/PfT5CzMR/
F4rbBVbP5Nj+6tA+5VNwyb5sTTQfGWScP+Tf+SW60vGEzApYEgbqCg8DkC/tjhv/DORJJvOAdUWa
s9dfpMooMyNMA/R5sqVuq2PuRVfAGdNX6ux9fAzM6TXrGz3mr0ioOSWAGfnElc9XvN2a17w0XBaz
Ct1Ly+Ri+Ddrt7EoQm4qG2Uo1S7PhAiCrJ5BnwLMH63OxqvJGfSyIye1sNbc24kyCQzfBw8ELQwi
o7qlUy/ydv5lm/ILFjbLbiEBIPuq4d0ggB2kKF/Cy3hefvp66pvZPjb7aF6PiL5XjGV477DBNDaP
si+ufMmLKOIlhm2VFt8WDMOguGCUnEVzJnxAJDjX8PhVzEBmTZ0yWZ2tI6tumc6wB6CbTw4Gza91
drNOrAniUP+ryMJv9A7FBo+lYkin/54X5i5ScnCXVd64jGH2BedvD7INGKrtBsqJkgqr6purhv+S
xLZ8iOxh7j6gA4AKI5DI8DleGgzr6QHzkE9+O8c9R+zOWtvGhFZqaYobK9bXnRAVaZxluBuOSsLd
J/ZrwR51Pm7jsN1oeYCgySReY51sU4xAZDYlSimv3ORWMyJxh5Bczzz8tBY30NcYn03HJyjhKtvs
XwHK/2d1zk1qP1le31IweW6mFnmDwVJfACUvAy7GX83Zpgu9HCwyTnBiE3IQSadSgnREBsXYzVJR
g0E69Dyv22okmtZ96Mk1zYbJ2iVoWUx3WGI6TbOzFMJoQC9DCyFbl6LB9hJ9JOjSW5DDAG5XM4if
uYL0Tr3ItexUfTKo0l80Z4Zic9bo79e+9I9cErKyWDJgSh9rBF/gT1jwlTU+MuXfYk5WRME6VxiQ
rzlM3D2U+t7q6IUNwFgAltX0r3ysnBAgm/lDJbTibZkDJImmznFEQbGhtXsHHwKVpS8EwcLLcn8V
dUSOhn1dqw2fjsxJQ+Gxi5+dNQDPQku0hheybhxHE1BDfCGyWIiv44W6ehUcpZPua9hMYphr1mS9
PsIoW5BxkxcG13HdC5GLhSPVwo1CVz6rEWnkcY+xZYGxXitbLWAouLyS/pncDT2UHE859Y09dMuI
9PZwg3tN/XBQ8nwfPqRp5uLPNi3vII0KYo+TFl9gm3nbweRc/UMTYy3b+iKMIGfjcHJkaD6tdZmH
eCGNTPZ5Qf2V3gsixL1N5CWNU6OUqDkvgDTVa2aKKigGSFAqsrnmMevEBkkZu/QEsam/uATPZGPy
2S5peuhqtiqGDnGcjt2T2WHF77bAvonVaFnM82sfKmCxQLgdFiGmMX9h4zTJpewm07S5YkYMuMXa
+6uf5OutbCvMUxdt02YNJ5DfeUWv9PgcNovTFq4D3dJiPcI7A+VQZcRiJyhlfT0fmsOM9dr7BvkR
xdcL1+v/tWqm3bS9fHcqIWAQCmzh1RSPpVgZpND+UZFvC0dLUivSiXczX1KEqONUbJlXb0llC7Hr
JAADi/C1mMQPdPyqZLK7BPBit9JlTHIAhWUmzHug4g55AxlpaLbXxLTX47Hk9JgWBc8t8I1ajNX9
qiMdHHs2cEWsmJI/y8ynUscq60iT8AajbFnklJeFV3au7FCL1ry8TrUpVDEnHvBh547We9xfGaGx
PHj7eJS+K+hu1H4Hbf9Gbx7eIwUo0znscGSuQFhXrAcCc2/7EOnSEe8dO59ObeUeY8kG9fnGArK4
RBIWA45WgKW8vCx0V+AYng0ZvJwFQchepuMxe4+9dss8AZFGTgSFOLEQgxwRj83h2KC/m5PvHnQ1
yfhBsRNNuZ/kKLlMmiubDJnFgGS9D1nSDa4L1LlBjHL8WOetZn5h1/iuCC0l94Jvxpvx/SDdumct
D4lPp91ojZ8+jaoecGCh+G1Fwi7jNeEjxbCVUjOULwQtOGR0r2ZNgsCjyulzVJ8OyY2+7XK3ZY6s
9km+OlQBlQF5KW5xgIIY0tGMzKaf9NTV+wt8Z8EJKuzgTX0kEvauvOLAtoE33k3tC19ThRir+iZn
a0N3jobb+JSpMKIWXEk2z68J0AQABATVcFlU6h0K2kG6+LgA1UxK0he71/HFUXWnN5w3x7An9I9r
jUa7oDSUvEXPMzfVe9ocqyhfqBko1o7DVYaAUhVIlwk8ojjGlcTzi5q7nVYtPSKhIOlikZ8I3EVD
CX7F0Cu3B6B0AH247uNXf5E0raerqD37Qm5jWv2eY7zTtTdLP9ukjC98s9vMmeSl6ghvkp9KRApx
a+bjHHCDj9j+DPG/D2oCySKcO0XCHT7B+DSPsxTDVO1jwhobAxRFTzf9Nt08/aGepulZBLbYE3+z
EJrBZQbK2lJ+gdfuKr1nEOfzEe2gtdwlFgHG4XR7PkEMPf2HPCinQDxQ+gcpdMx75eI1dE3FSxrx
dtz8wuPu1KyR6LobeaB+C5/epM4BZuEZlFi/AQUCi/DHx/jBv4MU8Kw1usEesnEYwF2F1nNNzmBC
fRr4rgd7yWI/xNN3gHVKCWzIIQEwtDI1oHK2gtYquigX/G1IO2gcriYruf7nFno4XsM99GgIs1yo
YcIgeR/ZSLZqwP3xjX+i8S6xo2nzYuXJt3BPcrnD37cJ1mLXVzK82eCdqez1vQlFMVEOTlz9c4V/
Fvd6XGcQB6Ou5XrxX7jdhg0RBk81ZDEAeATMAh0n6iUIFl/+DX8kGwkcwKAxQORXJqV9sq1yiZpW
fb+eqoUFuZq2n58oDBUM7Il1cTAMP7gYb6v0Fsbfvmgxa6bGsGFb6RZ+qKUdQ0bl3yZb9XRmRcf0
nkxJMQxf0fSZf233P0UtJ1EcW9w2JZkNLWCPSomHxQYIHED1W0ABjlW9mUvuYYWyqg28iq5SZBTb
TUSpi9mf2aW7BrYCOuwTInWPMQjCVGmKzoGl4XQzMM0P56ZqPc1eVM0hQqkHNolIVhw+LSsE+iE8
qwBgkeBcetYX31wjvsnO3gI3sKW2GpCldeLlXWPJxSldT+SHk9d8VlKGcMj0NP/9L4YHoMbwVgNI
0aHa/ypIesSL7JK/08RwgcOqxO0mJVkF6bjDNg/dhU5Fi/VmX8rst2acwpwy7/B48SApIQDw0YgE
n3QAQu1YNmmlYS98jBNzs7WmzYO9h/wefTUxEbClglhJxXbc3W7npvPVU+4H0l74HmyWrePX5huG
/Ofm8iZ+vDhgtduQhhCa3T3xMr33hVnnsASRG+i5o55iA+p2K9zuTXf+woOHVe9CTKE7Da0jCEWT
Bmx6ALtqGUpspvwxPHOcFWzPUmMIfrdrOsJ1wshRxaGXjAAE8s8eSCVAfAt77l1gJYum3FD8E7eS
/eV7M4C67AH14Lz+F2Uaz4yyaWrqdOapfkh9JPfocGoHPUITWr94IwhXiKHDRkEdQ0yz06X0b5kq
+AXDakGT14BLJA2LttP2J1GxUmg5Yf99+5/eq4818a6M3qWQIkJb45/6bI9EF9tWBDJnnTSOnQpP
/K4QRDz0KtyHLWfqEdGD5eFAOkC4mfXhK4YLC64hryNJ5h9WIkB8riPKdov6Jr+cD3soFoypHCrP
sqvQxRnvpjUywaDbjXI61EyogaVETndHoEj3fcl0w4undHnsTfNDVV0e4GK03mvGBl3DH4Ro2h00
ib8tfJEdOP1wykgUx//gpp5of1A6BbInvwLNRGty2KiULFhmT/U+FzVE4TIGvDVrwBaujEu3SGIC
6R8NQrARYpez8R+2lPHo28M+PoSfteZgxj1uNdQwvbHv16+GkCDY7iOHRrMU01qOEovEs0f0bLBc
CE7mPEGOW/wGZalqFHXeL73+EPBtXLwFY4PHzyQq6QRw5ECBcURaPs6yErgnO0VX0D7bKVfSPKM7
z2/314IhJ3PRzCeM16pxJMuXR0d+K/79yTvyi3HTkc55Zac0myGPtMm58q3kVX8DONXLf6+kx/qC
S+JwhtkDYXkOyJKnn0UmnnI9wQ4CPoXxLZUHW+KNS/y9t5CerL00dEaucn1eoNIxxw1Wx/TeDkVi
5psZM+CpQy/4XkVVUzBysLBJ0uRoxsbJry73H60xK4AFeaZ0bj6xwelOvYUeM7hxtbYHiWSG+pVz
GJCqG1V/2zrsBMeM/aZiPK6lkXxt6/Lba0C4nneav/+G4UhxH3oDd0xD5boLpP96L8KS3hNLKeCu
llEqvloigP1xp3wDkPYmQGXze1CIyZ4QwY1m6qdllBK75ZKO0gLl//NnIuRyndNutFviBoubMS7W
gM9dA852YT/nAn8G6Ogb9VdUudr58xmPr2HJivvSIiD+WEDrNH7WM1AQ+nWw/eRVi+B7wD9kqCE+
PSf+TqYyouPLamSTViWm0bLfQW3VvkKn9hDRv7dgTht+V1I57pteTlNNyLa8xzWJRPAS83xDp1Hv
e1eG7UeIsyqE87pDUzEIMqKKTyh4EwU7N2myRF1gpx9apWG3M1ZNbLUs7mqjOjoEMithEiNPW+1m
l2NnWbp2k0mM6N1vzPlOHJfSUEZHkSih424ZQWrVm+tynVMuuLwQqBy7PeHPdItyPEUrWDyz6zuG
dBhXlD8SdgAnQghlP2voIDdu+jsM579JnWuLmWptrRJmxNcwu21VtHRqa3v7W3TIvumTrapI9Itk
J6rYB4MM+n/I6mzXNngRNCLDEDCGNpgcpdySXSxt7xVFZEpBU8205I+tRsalXPHpna9aHFbSLEEO
2kcmpG6m0xxWKudmVgy18NI6iJQFehM1XR1orxVKtCduS1k2ZeWxX+cVhKdLBRMa/LRXYwjFbzfy
nOCG/FfdqdGX9MzXpCfzhoZT05bJXzc0VMCDCoi/NR4h/rq8rZhvvogxaleK1IrZ3DxPFbrH3GKa
GmhYXuK/jmKoL9aHMi4K8Dpij8J8c59XMy1BSKv7U4Qb7lvdX9/rY0AAug1a+c7A1FionWRR6mz+
ShH2fFphrbBtlxhjTFj4XASBTTRRsETQwYxH1APDH1vng56R+2M66f35P2mdqTiLCMUgpf84vScW
ywbR7BKh8PDJsndyrTM6cXV3Oppd/3yCFhav8KjQbkxIxTKkODQS182ix18Rwso3ltyJhQvhlb96
jzdeh32RtS7fHXHbyCtassu6e6ugPA+PemfQWPNLdahQCVktiHHnvD75IcLRQDnwqBICKAYX6BNo
1G5xabCcypVEkNrMn8FDFdqhpaD7NkdOlnoo/AL4aEnsT/GaUjGpaSWMe+hVi7+CMyXn9Pjp/Ziw
36fsqGE2/tQlRx9mam5FMm4WXTkJGtUKbFrU8E1wMbP9kNJLeAWIMkbYfZO4SUpmK8l6VV80ekJQ
TqjlW/O7kLjvN4GYrxN9QOEX/6I349OMj8kibWMkqajjMN4lmOOkkci6FJZXyd7M+6V5p8u34eZ/
fUghxecvWzbm3dG+sI55MzSwwKTgj/E34WAwGhU0xqEs1Co0RbjchVQvgPW8Hxgworujd2WLp/TW
uH7Frg8q8j3m6GIysXqY/jSodu0O4w8DhCDpOCUy19hL7RsrQXBp1mIbEhgKtXvC8J8UHVfRLrds
Kl9NKfLxnzAgGS4lI99DdQ7o5ydjCrc6rQQ2lrFvsDPYfmcP2XyxF7QFPetwhjcsBsjB9nSxutz5
9P6v6SuAwpIyMug8STvo4WD3RBLWq7JGcnBf5zdsKCnl6N5Y1BV1nFniQYjD6zHw1kj8wGmgGx3I
6yZPeP+EndRDgT58hEgr1WZvppXFeT5Rq6vFNUpV+kjYdykgik+qVviOlYTK7ICe2BfRi7onCScE
QmS2Sx0Cd6hXPSJRHDNprPRmB/2c6BZmrQSSUuw/RlP366CBvFORooDLO11yw3gKhM7OgT020l1N
jIkqNRInT1rE6FmgNVGS8jDx8Jba08KjMsQY+63ywJ6lh0UTPXr5CSeBvl8YJlEU2SJNRdtIuHUq
XeeGIoQ5Jm7JjKchgJ6EWUM6pUuJtqja9P+ARIp7rfWT6B0WaEu1zqnWaPjVjHyDvJz67YG5xCNi
7o5nUOSVINlR0x820xIHMAc7HNhD/OOs5yRGbfdCk++eOM9JTSvnLClft4J4qlnil9WXCkI+DvJQ
RnFdPqPOa0sun0Lph8qVHTgNiKXnVpRMYn2j43lCOcKdNADjf8RogeYsHipZ1SEQRIFnUMiLN5ja
WAKYgjkNzevN0VkN/vH/vB7ZJ3V/X8cX/crwbel7dAcYyNK6xzoq+BqMRN6FHj+AOB0C7R4iIkI/
X29wPA3IjefOr3DTsQ8zMVe+yg65KjAcbSX+Xh0MPCfdhwxnkj1ciuFlIX3Y3opDrj6z4ICSUXj9
gRA1JEEGrg6625EnvX1bccLiEq2UMIcdcUfhwzInuH9vVBqoponixRPhlPeXmNBn717YuFN/BLw6
rjMmCuG3RwxfiMuNzllkoqCNkqNM9yUmPhzzVupSOxwGwFmeHq2ZzzWrZ6RIbBwxVbsBL4zD+z1X
fasDyxzPJqeufcTGAXT058hsm60kVBLEewBhvytOTlc5jgVtfexGK3GK9zkff6EDCKOiM+0Gj/Xf
pXx43HC0j5kOHmVN0CT802ACXo56lJ/+Fvr5qd4g9Dp2YF7llQbYZxygcVTl4SN4Df2XONl3cIb9
hXDGr0WR+YJGs+3So7LaU9cGS7cDtui3usAHwMJf3RtwxFu2ygH0CHfjX9rEjCPyLEuL0nfRPrm2
P8axWyCfMQ5BpDp2rSJngmKG0WsgzFrOEEaDPocfFzNefxHV+20oSTQpFViY8kdsUVgDsLqzbQhN
jLFvFk0Nw+w+/MY2MjU5JaIsi8NuIAQhgedHP0mQu2KjrTX9+C6Y4nXtTjxuU5qBIBXyoGArXvSB
EAldKYyujbvl7EfIf/hvB/PH0iD7K1G7zDjxeFx0bGnj5sqqJ4r72guFQ7Bxmx7QvN0VSJ6Pacwp
HPPHG722wM6LtPqOA9FuB00Pu3Fy17cmD6jy/sz30oGnPYhDKNoDXH0NcUlCXwcI/tZHbuxQLrpM
iAsgX0aS/JcTu5yhElvMaElsXUu0w/waVprV5n4RghElBpFjTz5DGgLYSMVTWJnqPc+8vILelPT+
G/ESsgbr8SlRDS+O7iGpA0Cvb8Cg28g86xs345qriXAlgczRtXcUXwNfPBNw+ICUVIVcw6PjCnyX
IHtYwId/XLL3pYYbkirmS+57qT5OYs7qRWqr9egIxT3aywe+/B8AAq9L94eXU7SeGJoZYGSBDkAK
hXvBA4QESdu1Km2kXl4EhO1A+7zur5s98+OFee80SmmHjvxPe/NvUmeH0EKJkN8ajqlyQbt9g8Sn
KQ9GZenKXapsqYldxXdauw5daa1lDBFKay0Ra1zPyDoXKHObK9dfIoH205QMRDtcs0zwD3Hbmc3A
MRhdlL0Jb/ddKjkuKbBnJ4iUfHsCjTXWGlO8l/BHIFWOm1VDXlH1fAr3iKZo+VRgS5ao3t5/X7VR
vqR8gLOOE7Eafrv52nUSCniRNIh3jT4V5WkRbRBw2ujCSJmyZngTkhkGjQce8r6J3zFrOjoe0YSG
A1B4mZDzxKExvzOsQmIZgSjKy/eDbS2EyYc+M+2ZCBGbd6B7m/M43s6mYT5U22gqUbXyGy6b693C
a6pJ+F8YsA4/CQCkAsXUbcv5MgHFPVIcn7j24ENNQCpOkAEvogQVaNEzslEy0B+NbdoQ8vvkDq4b
PeoWg1ksSrBHzQUFWzPN9zVsCL8Vt7DhsYV1Mrj4jy3BtYdkIfo0wme9xh8gyGDpN/EnPSaeF4/f
xsMkQQTT6MfYRb4MkLeqDpFMpncOfRRf45GVeeulblt3eK6ndkhyryuFf6IaM/Ev0LT+jwtC1bfU
GBxBit25GDWbfzzJiczir44hCqa4OvwELX1BlAOuVQc3r9INB6HGIHSqciqoGAe/PR1QQ3XMQAh3
4UJD1K7LG6ObFfMx0aW+tc2gdFYvndmY7DCVCeW+YBPYQkP9ywG5pgS9FToKnxgWZd3NQ+tuoIrl
1fGgS8ZdBgkIt9VbNnPIsSrFB3HBcg+eT6W8IZlVweMIcG4tKcHkbKgOnpwktg3DPpaWgreF5Cwi
1+TvfwVWfGgHUubcXFcuS9+bZLOB5iUMGFaPC+nEYVgXGx7NcCQNXl85gRxSCm+UWC0R5yFYjI6a
Q1svKt8dYp6VoW3/yhltX7dWrVbjxJEUdVruXWtVpOm7nXQZiFlfcVla/FWaRhKVvw7ox99iQoFq
1XHFDoewoLo3KqxQXa1xYBddoPye5v9VKCid021TOrAKy1ANYg3mfPEVJg/FAQXuKDuAjtx17RHN
h9BlL91fKgXd4trBc87i0pDSqiMU9mWnffZy0wOXIs/YGOV+rixn1yR6aFnj1oWnvjD7xwN87tlN
LWxHAzqDRdOmC7zS1/XZfUGHTS/m6ylMz5wDcrq6jTube6wHNbE1sHM3KwQkibWOgW61BWGen/aw
kvCnVUh/6LnubWDBRmYnCxAgINwfREQBY8B2Kss2y/IJ+mTscphkfROBLx4+SUibKrqBIAHsiV6J
fVrLfRlopFqYUsTn21iW2E8zEWCBdtpQITXUxCfW42y4hvZ5JIjFFffdxG/zg8PfK+J1xh02pkOP
YbAGZrmZD/+6nbTO9fj6jXNXPlbqduQQt0eVK6ku5gCmXt3C8uaWgi3jy0x6b5+b7Do37YHf3buI
QuVa7T+hjMkhQCA+TasimgJwinoeTQOST23WF/gqrKb0rAwFXf94sJT3i0sNeNVqvI0E/vyrhRat
e2xL44dmKXe7IjmWiXU95ilVaa28z8OMFjDzN1jpICbLaiYhyWonKMgPLBr4lcc6hSB2ypL6NMpc
SpOmJXlPhTRVR+6k5MFloxSysSNMejtqm8TB49io9/8r5lzJa8rP4RrsLAgyAv82cQ2fX+HhCV5M
Jr6YsI4Gz1mzfxicM/zZWgB5skxCKFSOvQXEIm+jfctAeskuPM7+kMEgMxw8W54jqvzm3AM2FF0j
KRK9TYBHvZo8NSrcT1eZ9/OCYQfyO8ipWiI0+pubiU2cRImzc9CfQc6Vf3x68Z5VdSi+vRL9doXZ
tNNfWa+ap9t9EYWA4t51dgJifVV/TM+OBCg6rZS9Gqa2ZFoABaaSMzCvqPgSNJxfB4rklB/CQOI0
/H7V6MOr3sCoyVGATVTlHy/+HxPfalKTWaouR5Kmh5R9K7lXv/wUXOwDPX92bgEhAY1ZPSTa/WGY
PYa0XmYaXvWGEQC9j4kr7oEC6luQUEzOu6dX350VgDVbKh0hjb4w9N7qcNR4P1pKqEYq58nA23il
H6nKMm1UvZTE+OCbJKWE7WQ3Pjk3iw8dNK7UHycHhQwyHMmBALHh4dHOqjbyVDB2rD1uW/ps0i2J
uPMoZ86u7cS7GRVenZkn/bXjdfUyc/Wzin2RFWpG4KF5LT5lqFtvRZ6ZtAJJexI4DlAGff0m8XOw
XgKfuBCHvUjGfDF9ShCjd0fAoajySufLtHxnBs0DP9b7xgXKn15e0rA/euj0GI3a8LoNSgKVVXJ/
tOvP61oK2jVP1Ka3KdTZAvpmKEM3bKPhQolITNxERGvLIXq5DWsleJDb1tpfy2egl1UIwaJVwm0X
c0VxatqLiQSVmvcVV7nsoTzLMq+L+QYH7wn58CxAr1YO1cRjdc/gaqkrMts7FgtwinTbCEj/p+r1
ZHR2J1bqx46eIjROMrsZh0poSrhVXGy6+rSu+LiygAbgqJGQ8LUFxi4OFUQ41IRR4vNfxBBCRb/B
tqO6p1QJnb64vmJwd0gLoACiDjdjWh6AXRdeT+f7UkFOFbwpsZvT23iW39bCPU952USesSn1D28C
6Zrr6xkUhsackesDPdVPs++orfntMSM/Ot6bGkxGdyyljSLWuAqshVZf68TwM11Ug3+pKvYnKTII
7UEjlJr8+hhas9mmiIxjlbuKS7pJoMolAZfeYdntvhTI6MDhFALgtkogydedpKt3L7dSEdI5cnyo
bkDoUEOGL5PhLvIkS2YQ7wC/mqwmm6ZXwwI3B0av51Ag47SjMYvo9q5pRKmjeyC7GXJbRWeMh/Nq
YAvNDbsZ7jAtYg0d+ICCE+0Y/uNONxOKAmmazuft9t1GE0PKzJsejadbpFhQOpDVkZ8n8eXg28RK
BYzlRY1YJYYH7eW6bCVk6N9NhKmMf2qwNAd47BfVVnak8u3/FY+VbxCghYNbZnC8y6vnIjvXTuG8
lxtv77trNDomrhMKUcdn6hUVEgsnUP+WM8LJI0ufk1ZAQg1E2+7hdM8IqskY7D4XB/PKOmCH0lon
5gbB0AKMiDll/xoj9/dAoPNa4dneodSGFL7XfxEKyJJRPLA7osq2gdClBDCZucoteVekswK9Yqd6
1cy9K3fCNTw6lCGcXD8Imcz7C9fOzhsn0ZJsRF1ue89iZqGw+ePhOnuJ4FY5t8E/aDSyWEnklZYV
bWxnmsmfpkk/F9a6H8MzUGRVbqvdLKPtV1wPLEQzR1ZuBkD69W2ZELrApvTkws76QXJLno/1jwCT
u9p9KOIrxyk+Kc8PlAjg05FNt9AKB/F68QdVHDcLscuuuqSOEwq2u3pA2MeKNrWxEBmeNeRWAfHs
qncB4obNR/Ciep/bej1MvU+gvun7N+RZQmBQXfzy9TGY3Szg4jYGtjnkxNrvjVq7PzoVXPLlj++x
0WeiCdcd02hGsW4Puht5QOEdw7E0GihzCA0zUmCihgcA0dNjzxUMRjWqnakyTWdFTmXzOBaqkTop
mfo2oIGSsw8Mw4TefraD+She9T9kkF+kb4WxofWfoK8RcVlDwr2y4ddg64mObKkP/65xQdZwlAnv
0pG2ZRUQ45RibUTOyIkx/HDwvcGgv8jkq3CVUyREj9KlLx7BAYWdNBJhCeQMtyDTIlUcdqJFLSjI
qwKcBrYVEIlkijjOACsLThD7Hze0OlI45uoVRv3PsiJ+8YD2NI6KTPJl2US7TWXcTH0K8vG02gJm
380z97JumoF+ro3md+fUlD1kb2VwMrc4yckvGVI8LDznsb+IKgofABb0An5ydZei5FvX2+K6pg0J
qpRyi0nmaRa2cxHWeoytqCWx3dRB/pjdnWBtcP4QmNQX9FqkWY4KrfoCjyX3dfxhNCeX8nNO7QCv
suigjgqR9lvfMEdGfVGVukDAkIOPcmg/92yBp+DcCE9K5Kz3tPlv4n+iQSYnqLjEiT0rKcS3GTgu
kkdqgKCE9FVEyC5b8o1qf1QQibCim4FnwPnVZqUqiNclgRKO02z7+SphCVBENg517J35PewUYBCM
XfS6Hb0Acz2w5Gl93DFKi+EGandbqFDxjpYkvV7WwoXJ26BzwfTqF9VlgKTpzRny64wly7+iqR0x
2RPcfze1y5wbJWIcPCYiP3UYByzbQyb+ud4mecyi/2MkqIhgGbLZ0QutFa/RnCPYWRcba4rzUdhz
d71wzg2XSDEGV5qsu6rMiUa3cyQlXHQV3avpI9ROhPLKJ9k/mZY99ru3lqbbiTdcOZw7LuiIh0d1
oDx2uZRpOfwGfZCnoB9q73WB4sqj384lZOIh+nEBEeZSNsVTRSRRfwD3mrV4MdgayEYkpVD97uOC
1X6Ou4tObhIo70FXw+sgwLJTIYfXFP1n1HmX64fJqqIAxxPqAiFIubR6azp4gTXeyoR/O0BNaqcj
UJJH2Pb5ccZpzGzUWmkkp+kS8TNoCpxJ/RtdiPMSQdnqMDX9w7Lz9kM89NKhFaAeYMzSIbg09w/f
tJ76CrUo1J9r1P3oHPhl/EpJeYFwF5ojVxN5i64OFbMGgBWrEzyN0nZ5nicoYnc6Iqvi+iJfrWx5
rXE3Bb/2vqa9gDgSjDdonTZ29NhDpAdKhOYNJI01N4inSbCF8Vanqcm1wzAU042GSPRgkglpgNFH
tUjI89LPlzcsZ6gEyJJoUG369yopQWdXwq6rjSGKH0vHCMiMAGz0YmByOyDmILUKbCRTDChr0+Fr
JLusmDGsz26pa+PD8LYaILa5SXvH3laoDi2PsFof/z/xZ2OEP8i0LM5j5R1viQP26+aRXmTwv+lC
ZgcPdozDMYW6uun+vgdmpebNmOmSQe60odZYsGEvDFB/L8YaumXjvH4gnVpMWr0CPJM7TLkQ92Sm
WLak0hYbPiWrMHTJLjMwAyePHs6vdkfJ3AAOUtUd+QRLDudbEDHHxjsQHKD7gf9ZP5K7qOtFC4qy
tMAfw9LIlPKCx1X4l46IeGFqmZ+iG8mvjY6SLnEtndKgvBlds8aoyyivopOOmpLjHy1AmHv4DKhP
8k94PeJTyPwfCh5SBYh9tBMBIWpQ1ymf8Ls3nb25TLCk4/FfTP+YLdWe+UNuhf5fN35MdsRrS+5j
6AsQElppFZYlBo95xwRQeNdF29WBeSS2DG9BJFCIaiKdjNTl42XrJgqeqf6HXceG3DhEpV/tvWV0
G17c+9/P13omKjh9uEtek9oyNJ4hQWjTwuRKF84K5cV1NOqtWyytsSWmfWpEAZr112O+ulvzcKx2
izHi8ZjCRE3W5hbE+TYTODz07nkfith3MjHzwpOHEtrxBk5ECyNyfDs7WZhtTSDI2lSewB36Zd5/
NZ1g0ueuCUI2HuL4Ckyc5whxNBMvd165az6QjZPOr9X7uELv1ZX4PTrOOYdZFbbxfRovmDk/p/Wt
GEC3yUOTb2SFjBTIesrbwAjdqQG9/f1B82al4JALNb0OCVZ4mQ3msMOfl+2Gfzcupk/p7v/r5YjL
mf6LbecmdbBGxC8xef/RS/GPHCGcYObeHUydTNbhAfSWmBf2awrtaOnS13uJmovFTJH2osH/kgWJ
VTZXH1jvXpDW6aBqJKc4x6HEpuoaJwMnEOzd+9MNe672gNRkQdse7IbrzoDv3KxT0USvBy0bziOd
MwSqF8SemLfO0kiaXRl9Pz62Qb+hwPcFFktYr6hLMngLwL6DKkmNRsZfaUSLQPRAHb7MlqYtDg5u
iORGtuou7U9CGNFtdoxpjWoKkeDJ/m2AnfGBDaeJQs8WXvafh4UkZUoTaMjRuvYGjwhTMTrb8/Is
YCeupOvHgD20X9g6M86ykDsb9AZxqynBIPFDXCkdkJxGP+UXP+DS8wWiFCF7u39dkSokSMcksdY/
+0C2sXUuGHNOkec3xQLoiyosMJcFg+MnwdHrBtnYfbFm1rmRiABVShfdwcqnRIbR2XywYJBgbR8q
Zs9ZajrTI6RmUfEb2WFtcFaXBYurKmTvphaP3SH1SpgjNcB4LcDuyNsou8Wy+m6t3jZOnuNkpfth
/sOL0xUEwDnrL5+18zrxazeFa3uQb1oPhIw81T7Ze+HHKcRoCGIYLt8LQd3jEUqj072V4hFBor2a
LLZHwoe+MVFdsN7oG97Y1Ugks83U3vpmKqtbBaPOkuLMJN/+k6+bE4pl2a6j9z4Kom8AnV5pFGhT
UaZoCvRA1iJu28jHKozJ8v1/aS/XtilG6giRD42j/lTnfe/nRaVp06uFdPxvIcaV7JBS3GSCcGgW
ve8X+cpnXaDqU5IWX6DwYzL9N2h7RGkM8xTS0kAcxPN1Jow8WQygbNXayQoXZoFnunZN3vp7r3Bw
hfxJHDXn34gmGjcY2PZDWLX1B2duJT+m2peUnJnaoRR9liqNjypOhXInWJl0BqUuyU48V30xF5Gq
ZhFQp/DViLRYJ4zCkiSveNeKBwDg+6eZ2AfHcCwBMBtJOSWosvsMDWZy3J1r5HJuiyyGvijXQBJs
D6OMbdlMxl3CEzWnfNrW9ANs1LTPfcrcFhdMCgX6sNwzFjrX2t8kkqiFG/B+kyIEFyxt+I8oCLL3
Wjxn8ZaXtMleL9MGhoj2IED5E/rY8cl4aeP1TuWCsRt+aTsyhqkaUgjy1sTvKENP6ErMsv+EO6Gl
uJEgX7cnt4sSnXEWDZD6XuVJ9jZcNi87k+g4jKJFxhMHt16F/qXsR/xOckVyT5SJOVi4m9h/s+zp
q3n7/8+x9Rd4wCDr3Res1FYpO46dwJGQbD/2bLvo7visIo1bzk+Fera0+MXuIEai+Kh9bDWfavo/
K7CJYURBBDP0n/UzK1dK8GJP+Q4KyO14TNfrny5U8wztNmdFVriV6ljEbQy1GcZywUrM4PmfceMh
163ySxECpuMobUmtZshDFKFqsSzN6xcifgUKMLJvrwqpEk9FetV5gF6yHx3TT0eUL6LigtxtBgdj
DkQVo79LNx3M2WL4qVJP9PPT1pza8RWU5v6fZRvyI1xHZ+pCxY0ooB5eYACIjQQCf/EDYTBgLUBz
8V8qYMqynWn38ruFSTXlpApRmxb4JZq1Ps3bjp+kggFnhuYfEcv65sYEmForREPppZO+qdu5Gg9M
9y1DHElbap/zzzTCzyiCuOrFLwyN9b4P0a4oIa+6kwhsPLko44fB/cnvgT/KmpGAqOThi6hTqfmp
TCjX+gKAdohKS1trlsvG5FCfsAnc9bmeWhZd4yRlAjW77GKFBUQ/5whBo9eL3D38yaECz+pnri02
OLCjcX0GBBYxWVxGXxWwRgX8NentAb+mg/oB2tQRndcdpAc9l+LG08ROH4NOgnS7PZ2gSjjDg3E5
+iSIaAB7V5ohPGx7Xmn48KQZTZcpl8riA15CodsPOZj9JLXD32fKo8w1M0H1Vvzkig1NnQ1xZcwB
+7ds6cksAUe6foyipSK9LM3Pw/b4k37IF6ZiW2KLTp87A3Ls3NukLAOAqASYSZztNfGdNFlMTWia
9NjGuYyfLNxW8FE4GYNtVWs+2KxnjeAiXUUZsQId+GJVvQU3vfPxj0LJCxJ1GwmR84JrEpuT3VON
ASrTZTNBFXEnb6uoFfpsrllvjOEf4ZJK52279RrtcjcxvbGkjVlekbpWb8LS4fXxL0VuivlGrKAu
FTFt469etOyuoEUu1ggZpPvbnE4k/IN3foMQ74W9wWcU4IP2ED0fsUIdNBiIDoR5YiNkuXUUUSSZ
9zoB7o3WD+aF87ItJzu+ahqQYM+hznVbfPwVRZFMUfWpFQSNnTScEUq/UYM4DNOegmc320iYJYMf
VOUadWnxOkiD6Ge3toBGsHaeOKqAg0rhL43Xw56+CjQ019m0vEsqTTg5mIo9nm7uaZrrvKhHe1lW
GtNv5gtqfDO3vTP1cl/lfUc3VPTdhcFj6ehM0picH9nB9GASKcoo68AehfDnq/789gSfbbmFet9J
vzOcMbip+2M1Yv1NqBv1PAIKpaTTHIdQF6TFGyrsxjasbIUr1Nbb/9gIQHhPUsqeZS3l/Ymh+nZG
VfZ1rMpksFM29IDp3U7wkLI9ASg+Zc97MQdcdKVAEC9wmkaKT3WuYKBDO+Jv+yNKvOJNR+CgghRq
hybD7NvR5tAf6CEfITOumBP3RhDHDyP1FQGPtnkywJLYw1fsKAoU8ZwPlLwq2K8NBEUXCgupNuOA
fjF6UD8nquNzMKl4xTDkiDWd8QCOUuMRzQwq7zgoNh5G+EPGfIKT7a0xbdcCiplWlDXP1DXoDo5c
ZO5T2iJ524n66Tb4zlXpYjHwSwrTqmnm1iBMPfLGv8FFsqcoG+NyYaeOgWyN5V0Hsl3MiNvgKvoI
0GDQyyhEEyuQkhBRy0hNAckjoDvORp14pUMTh+P1XmswvDEUpWaCsnr5VKR7XS5jJTMH9JK9iT3d
I6b0rvHJDPu0ivD5JN4xeO1DidaGvMOMRTtYpInxhXkY+6IprtKGB0GOL8ZBEXlgZbZcFuGSo5Sb
h1vbxskjVwqCe93h4dl8xwAV6++q2PIfu9nkUZIkztL3r3yxV4+HhV1kqWLIRrx/Gv2SFwvyqYQ8
jTWWcz/Cc+mEMdxWu5yquS8QeA4ozW5I0qtU+IFuyB7L8itNCHRHMW0+Kr+Tmx6FkpIUH1KSXBWW
9+HD4yBrz7FvQfiR/1DCu92s+qk6Zu/4mfbEKLaD9EsX6kr4vxA426+nLmAdxoejQhRvYPwJXRWJ
OqQDI/oOt4jHWvjI860i49enymMS4wVgcnVky0v0KlS2E9auy4spRGedqb+wCfLNkd9eRKK6wlS+
ZXPNricfo1kQ+I1PUL3J7c7Bl1rNLIXXGOvWfCrbzmyuuudq5yzc0EvTPZ5cApPz7DyWdWs7BhXb
4ukk2NStaBeWov0AIj1LZmzcGuUsWkvPCjqlnF/b1Iz/KVqdIV9cMEiEi7Xb79bsgfNVDUU/p/4r
Q0WRGc9MtsTMT8DhazPOHP+4LeGAkT33mTWop3GO1a6B99ZwxtiINt1WCZr67X5JR9HozSHXAHwT
X2t9ReSQhZwY/oSCj8H2Q2oJo0JbXp3rCKNNRvIh9YvGdtKNL4/UUBQWfZppQL6GxnwRck7KheDX
2iBaJjaQadecoT/Fhxi9KKgyJ6TeatFavPS/ZTunujSNW7o8BtDftHlE9xjfbWigpaZtDefXLX2d
DJgFSOJAeGdXYpveJp1vRcfViXMtCf4JjVYqy4fwwGD0/9RKr9huPqR4fGkncKbbXeZlf06lpq1O
16N1ltyPLicVvpfryROxtepV0sEpuVFFqlPWI+kgZC/ZLHZB+hUzOH1m7A4cZRsnXN0LlBGZiIjq
F/Jz1UhbuC2WLwPYrcJL1WN1bXkYp9bXtBvR4IAy8ZG9wKlqAv1a9rpZrzI7NZDjhBQjdWEVxIlt
Dl/zn3fSdW3R6UvAgMwSNMSviHOy62MjKSNImm9GQhXey2EO7tMjly0laCICTSEK3VL3vkdItmUU
PtuK4W6atiFlNr2pFgo7DeGZ33P3CMLgqL5T6v6zEjJAGX5hKOawxnSfBic1Wg9JmBrtUjL7203m
EOXBrl0mV551F/A3yqakKOtLqcYPGL+B0CSR/mGrQxKASKKiRYC0TvPE8VvGmDwq3NXgLEeZAT3Y
iYSUbQR8QqhyTI/YrMWPhSVdBpNfELY1ZGaMGl3d8niXBgG21W2Cy4+/xo454FWPsAVjpToipMJm
CV382VIj4rLxgwX1Z2L0ELGE/apflDZTVcLW3Ojf28oTs0aH4k5n9uh/UnjSNmJZEJ7J1kHwx6Gd
kYsRTJAdKuFrmYLh1D8ZPmZ5aqp+jPKL3jzk2dOyVUXOxhVng1Kvtu8Yx51dXL0Gwl3u/eoQQLKD
MRPohriu1Jecdp7igwRXyNki0kxvzq3W5HFVQGiyHKcbTXoxj5sCi6/1x3VVS0szO0FfB6fDgpQX
bc/cGA8KrAIyA0IwYSKM3aTvt0wr+vfS8gJJrTvUEtbGH2vWFXYkeQ1ldZNvyWtcMHXN5QdmUFn0
EqIETtBEiq2hE7PLoDMxeM32D59MP9ip+TmMjssy+UhprjTBdysfQ3VPhWzBlzGrQHn1gDfJ/B9b
RinAwFQB1zx5VurX39obKtBY+yKp0CsMiAZf/WubfLRc1Hh9lgzCyCz79nZ3sjB+OvRwW9EKg6cs
qGFamSNfggbLR0lph6iiL2bhPUoUPaXzRMW02Bvqh3RQhBH6Z0Rs1lRYxiKDNcACPN2ISPKAQNyg
wvGFdXZvRdV4vDtmgiZ8zvW2UlOCJHjPFSeYI40u4kUfXvEdQX/X7HUwYeZMsfFYxRzkvsoHkjKK
PVGbadcLC9pBpAwNuHyCpRmJt16IssW9HL6qkUzLv0Li8koVH3s0qS69w4VtXl2jc+ZQG7F5x0zq
uuJ7OEiIfBJQB7p6k6XAWm3BvfmXyrCzz1llqvRnddh1S8/0aFY4HksPKgjaJQssRSwUz29Frw+B
GQwT8Ag+3igyVr6qZN03aPUG5MzEkg2J8+E8KJAAWLKsXflJfzSdt0QnCtGBg3vmf2P3VzIvqUM3
7TXmWxNqeJlutqz0z8/gsrrfO0TbJIp1c3m0r3LluTc63ASwqB21C+X0ivh5KnANj+T0cUr32+Gw
AtDNDHs8/Jtypj28w1Vrszk2TES61AD07iZOrYIVMLrzJvFJ8IGvLWpNDYLeytUfEo9rPKX2g314
zjTnCWW7xKv6jYPeS6sWUv8isltJEYqqrROElJDt2sJJzWCcifrZ5IPukH/aZDHPHtteszQ/CXTd
zcc8vIgKw0SFZ3yelmYICdlcvEJx6cVy+WREKzKhNF4LJeB3wpXrxEBL5sFBXmwLaje+tr9zlJD+
u6tOs658flGEL5TQM3TxXLwe3iocuJX4LlBFqqe782+aViFgxojOjzsCCtBnhs6vfhrXzZ1cTHKy
Bz8tR2aHtrA1LgLdG0ZCA/wIzw9ngQDUwQo2b5pUhdVT1dJV54P1O5F2mBtkRtRTg63rAEd3NaD3
J4catrhr4MTyDuhcHsw+ffCEiU6k07T0y1CLaSEGxmeRgjYJloF9anHFEvSvbUyZPR7UeN5LZ5Sv
A4MGa5i2k6MxJz/CQZurzpTta1vEtuPngHK4smQsDHDXgXc8Bqz0owps57O7BeyBoOqaGNFDfh0F
6NjTRrgQW/c5QNApkDBow6/ZWWC7HBYUP3HcSTGB1Z9eBiHPJTJZX5Q01IBie0CxW3SpTlxfQXCu
YalrRmb5Z57bUfBMsec5vZ6k6+4XW/1tyWR4H5WWdqppCW4Zw2E+swGwgEu8IweEK6sn4kNkUCXI
JMiQK8D/3v7E110E4is+akFOtKX9tF2/Kk/JLLZWOSrWEGIrw4guRxYjnWj3Om0f938sMHf5NPm1
dRHRi1DZAa6hW1H6HP0KyLr87V4ruu35vB/PWgILKX5NWCr2n5dPuHul9vP2Z5ll/dzlLa3xIZMN
na9gqqN1OGQ+FD2hG9t8sRJowjwzF1SNdWmwBpt/t11j/hHvOB1ePPlei/YXL/RV6isYtT+0tjmx
P3m5hj9KSsVC4KprH96ilAeb8DDA5cQtvT15CwMyDkPHK98xyrR7XeV79pZFUj6DqdK7LBlQMK6G
AgyiXKU8f7mdGemGHmY5yTmKVOb2pRwkxOfZHrJnah61EO1A44Tht1+NKX6ryhsFZ05hH9yHGs7+
UZVhPlj6JV/pw/E1rJyIhXuXIYBXZtQARlQAL8Cmzen5AKEKruBAZzT0mqEWWNcsxcBzttfEAr+K
iMfEa2ffTFzz5I5f/X+RyMpBg1zAV4Zh3XghcPBCwm62FwiX/TjH4uIWlldR7YzvpyLDMS1Vhkor
EorNwNhSBZ14EBK6keLcweoe74TDc7MqDV2huUwlI/FQvJWHcX+4hl4+kVKc/mXKRNRIX+gDKThJ
zn8tC/3CnAhXJ4bxAqZ56naXFntUb7rYXaCP9U8URS8rhvZJ7y+1uH9VxETWAv0/sKgfFe5Ytjl4
/f2EsF+mekcxsV9f744fGymwpqbeQ2g0toJxZskwJ/h7qTOc6ZzpbOurElhWEikFE/BuBQV27Q5s
3oSc+6WzsB9BrC2s2jhuFTr1/lHEYXBUXUIvpTr4rR31YR/gzkvtw6bjRyS89Al2cHuU3fC7b1RR
/Tq6/2FH4UVKaAljqrovwJ1DZHkNof3Oj0yupisq5z9uHTGJjyw1rPum89cFBPlZGYXrTPbH/Q2+
wKkDD9Uptj6q+8NdqQ7IbWFxLu/jE3UKemh9hTm/mD0ZTL7T07MDSDL3tUIZNKF/Ldzal+NT8kQ5
IyqzURcA0mTp9ECuQXjTbEIlbm45jko8V+pIHWSmYFS2yesRcsbApzKSRsn9pB/fjErhTMeUaF9x
5WeR7DbeWHylzBOSFHQAZ5jGNQqtDrZr6xEuuiAdo2Kjm57fAGlyOsrl70E9RgYGhAjuysWNTWzt
m3U1vqTX3PM6yRTtGtYUcdbtOJU9nrCBuQh/nkR0N9CG3eZEIH5aJjxA965SOjel4WXcBJgbkc1g
6ANg2XDB6dNgnKSE+le9/76zOxb/j0iNkAU2Wfri8hPjGM/5yBxeKsn2RXFkjrzYjkZG0ivys2Z3
luZrieVOLL/eIZPcfF3SO7wEsHzHmYXMF3iVwZ/f89HR8k3Mlw9/ef2pYbIozOx58NG9cogjtQ6g
8p9Cq7etyFrO2eUR/pwK879ki9jeW9sbR0hbcwkWzpoYT7E0Js8dRI5164UOZ0tEFsV/LLWje0CI
3h+UxG2ZRtdS+/YSRnUOX8JB20BuFdvNYF2gwoOmw6Dz48nG9DR6LOp6EobDrW+4m8AaqVpDNGYr
xvyBFS3TU5GV9rHobsbe5nRyqeg2ZfvmyeS2mFroKxYp5xRjDI0PARNzVTySdTeIibje85NFFEI+
P+wyOWOR029OsKbsD2BnpFM91/N4vmFe5t+LtCPuF0JnPy4X5AoA/idDKGc7SGrBDYvSZyvpy7CA
xN2oUJLgO+58Pz/uttMQHCikjc0KfGh3Or1qbv79R1cZoNpXrZUhAOErpe2F2w+ugHYw1jYecEKx
TvZlS95t0fOTwD8GniEb0MMDt7Mr29nfGssLRFpc2emOb9JHQZxkierjjvuzW6chnd0gaS26Ify+
AkFpkvc1k6uIKIniYelaMhg7i/5vw3Ucye05guWLKFH4nvHDub5Wrg6qWtiydQ9g+tuE+ECff8mm
jgUqvHeBsLI7uv6dcVKqD/Q7mWD55dGiuadgcdDT90dhbW2lUxSzOva1Di3g2hPr1KynbWer6gql
q+NjuhUHCaI4hilOtlDKY7o+Ctsd6NcK+qc6pIxOrYNjECGttiNLVtF9npAe8QmlKIcdVvwA6LiW
3Xkpi/LGa5H4CY3UXAwIlN/McPTdIJDM/q6yLEqvY9gMD+xOCJJlycPDHoRw1JM+0fDZnBYyXtiW
c9N5VRikUUyDptPxnWsqCEKMeCRbfI1WdK0Hne61vi+3HMrqZ9KGBC+lG85O0KdtMA20blxT14Zf
8hEZBf3AcOCVp2MJKOOZHkmgLxosBp+CKazW3UK/byFYGBttkhDQ17HhA+CcinWfVp9uXzXHGLT6
DGPDQPra9OR6P3MnDLoELyilDxmKPH3isGg9vY4UvKfjj9+16q2FAed+ULWFUpiicq+yuZ8O2P+k
N3fFqSiMlbZCuE0r1w+Z7PXYM6tHL/Yf6wFR1U5f3uOjMuFZtLHNzn9bo3VFIyAayeCF6s+zjAUb
NXsD6GkIO1CarMo6pCGuu7BKh/sZNydHCHXKkvWfwrpon2BRHhk+Ah3U/7lm3385rnA2WYeC3epx
1+oQiHutqnX4lwy9iSLACahX2VamtB9+jSLr5yOHFF7LBywZySHMvGGN6ERqBraQs4lPk+Baqw2m
G3ybmecshIyNLoDJnBnrWcyHZiWBub4inKYTgSQQhaUx40HCpvJ6ngCVmhJBi/7DovzF4nqqLlHX
BAmNum4RXc2BDFwrWA5zVlY4dOJYBWweg6Hm2ekBc3C7HIW8TGzF/f1bJA+JbhE2CyZnRa5vdNgK
zk6x3ufgVwjhW6XRKahuw+os5Rqc0i/UiGW2C6onqmrIxrky8Sr4dTxk15RBDS5HqsrOguCoPCCq
cDK+C19buhrDsuWVAlfW6XH7II8IGJScMWlbNnfFgSksT+WGjAvUd0OozfTH6DKZqcHh0MPDIeZU
0+bLiq2wBovoyk90iCacvO7CMzxbTa+8gH+QMljHsUX7xFH3J3x8Jmp3vxrMDxRPZUpvgwmYnMu6
k9EyN6mrOPyMOdHxe9/YtUadyvEmYpLVHZLThyAGd8iBIjfauVdKgJZVWJcjcnC7tw/cZIRI1At3
Kr0jbCSc8j8ZNspgsHILMmwy5n8NpVpoizWVv8osFpinPr4cxhoBrNZnx3AbqtFJifZ1sWpB5y5l
QBqOe1QLIeh+BU5wStEBeq29hi0Q/q6z1fF6aTGzkXeFXCj9z/lo5WGESY3LF3RTAjcP1I5Glnl4
+l2AoSm5pEYv+qXXtwN5Ht2Ewx94jxg2jspJGyPAgCsB4HTFK+KSLol/Rn3v0Xz1pqEJT1kTUb9s
fDRkxFStT8+45ENYPwr9S1Z8r2rdGNGq7raeGk+Y7g8tlLM55ZMwpb9h9PBR8pjByRCXB/801o6Q
GavBUvxGDL3wKFcXa+FA1ZFxDFTklchyIvGqHupQCzADYwpu+LQyMfF9VaZp1z9fE7y5lePc2Ug2
jOIp7n3AjNKKFiUPOWyd/jrAvYrRs+1E2QWLd3p8UFx06VzYXKH6mH/kYnpkd8XBgkWMG82IV4DE
NT0k6rAZxgEEn/6HJlt/Rj8MY/l5w99GuV5GaMV2eWuN7cDmDRNv9Of33VlWC1xGOkJJMHBsSitj
+eHWKgtRwYjHFWadenoSRvsjgo/94Zxq6F45/Gp2rytxFRittc6wfYR07SCnUS8TyXp+PP3W9nAa
RX62ABwlGbVTLHzkEERBuEJtwVbmZ35w3an0+NNwYvpTQgnsoSmVMlqL2waIKNMLUJfU8QE30u4m
mdPZGXs+ZKmBnVavVRBQRNxuv0RuEJXRwPbmrKeC0YReDk6gWRBLBXVDY8mNOj21dRs3BpyKcOMZ
KMEnPKKOoO7SNhzYvMKV4Zn8R0ZvPeMn/g5H9hzvriucrFAR+C89KW2bMLgDNorOpspix1WSvNGP
7IzRkvSQQd1/FTpppYDoX0e8HI7YBveV+b3CNXcp/wriP6pEhypXuvjz1nxW0UvWOerlIO94QsKY
3SJ+P3OGNRGQ5TYcMuPHoECI+YY/Nmu3UvlYrE/FpIgEAWnTLJ3Yj+w1hl8CW/lq3l3mbCv/s2D2
tbW02xERrSUdWqcCIkV5UN+Ot9O0TyEn/vTgHdlJHDDJ/2pGAXqIvNv8Z57P+3VSCIx32DevtkcK
MFLmyIn4PKD9Bg/brOdIhYsgaJ/lpE/bdZLOh6v9K8UnZ3iy27P5+7AFTiady7aQb+dCaOLd9pkD
4itni5XUUcW+XoSLTGueUb5Vm0L37bM3bAJH1exwuEtT8WU/6orf6MIIIxwAEr2169E6Hc99FpXk
hKsYG4EqJGD+JOyvcBZ2tX3TWe94G+IcF9tQ6A/Zv1mKOsXdpCPV1hS49J9R0iznpJSlkRjljd3Y
ZIJDZMFyVAZ78Lhw5cx1aXCrRL44e9WFP1FCzwC7jz3zkU+GyC5BYJBvRV3A6A7CLMLuXyb2pjQh
NCawmy8gtSmdZyGAIO8cI2Tj1gOLLe/Cjqe9yikuqFqIGhuzvmQo+BNNFrz1/kKCfC+OJo+AUEUT
QKqnUqJdblbYYQ2tQRAzL0SDD8EKqz2X3RETMYmdsf+AAvQrT73ndnvk/IQfGW7lqAg78P2Wd0wG
iSIlnpUIJLQad0nsZHpX/O9RfhkffwEns12KAZcrN3YfNzz5pqMXAO2w14Oovd6uXkLJgrrdKWcz
LEjGZLhaPiWzIxumk/x4en6Oa8yWFPqxof5x6CHYpcN3ecOE5yGDYIosJoQ6CHvhN9Cd/sjeScJn
WP9388cQWewcLr0fA4sYYutv+Zd1PTr9dKlhgBU2SabcXg4FopMkmlQEb/F4Vck7BnU0hQTAdEIb
4qunNOBcJ9YRw/EF+pGnox/tK+aIP4ZJKmZ9AhDeYFJbdtUUA3ElUAJMmSgUFGOgH7qjt0KL4/+O
+EG0IjllFn/DJPQ8xse3z09h01pDpeHqXZjbp2C9Jl16LQMnWNEZUTctIGXOYn4V3VaJXLGn9mtM
aROPLtMRzzTv2wQ42Xtw6bsEwMpMCzJo8GtO1n0ZRMElJ8AkiUbBLpkW+iFYi53u+R+DLf8fecrq
mLbUOK+daj9z2sqe98nEuHPb+j26BMZaDkUVtr9zaZXIaJL8W6uXfNfhllb5GZCYgoSvzGllU+K2
eSb0XwtpxyXgZr96NYDqox+WF2r9TKcXGGmELDw/PwyKNyjxuynl2G1dxnTzGNr6ppv/2G+OP3RO
sEiV5CFzaiZvePl91ZIZ2keWH77EnikbqXKvuDcGgXThiYnVtbVDzevlPj7FJTk1BtvN9D+AK36D
ANMIGGhYG2z9hPlEN7HrqjjUlSmX9MXcRRmRvWR/2Oz4Sn/ewhlavzg66fx7fO+muvsRo5XbZnBm
cd4NwqclxHap1z4b4Cflt+zxs5OpMvZ8iImtCXa7pQaUCMY2cyRRgctBcwcyDITt2BnwybRi4bVk
afHFFKdKF5HfdaPghtb/a/l/Kx85mThK+ZdBOy0ca++T/50B/zOLgdlfE+fHBg7pxDzdU6Tef0L7
vnGFZe5T5zpX2nlqrne0qVAwNK3NGcxCTENnQu3dNhNW63fCoNyXdiN/Qsu7eHT6JHnlG5Xf7iGv
4JQ7xqhZTA0bJeE/6wpU6H1hnP20rU6WdmbCiSdgsm9EWufIua1zY38xa5RrzaXt6x3e7Zme/t80
bT8GvdP7q4+23gtjdoGW0ZvSaRtHNWYEIdeKvBlKE9w0+KRqKlKBnaqKPdwCFSu84ygzHezhllhv
cSpF5iTs1QzeE7+CGnL07RTBQ3LL4pcoDBwxMXLXViJ0C3SNM0m0i8oelvXjy0g8owuJUj0O9nhA
zDD3YbB2ObQ71R/gXzrGVUmTs+w4SifwbgLqbasYXTeeW5cWRcieqp3LFbOYtbsIhCg79HPB7BRE
S25tVO++CTAFxQFYNjjoNMAvieLNSp5/iGIv9HWzLShaKqd1wEfWoK5qMuzqbRbqcQ6rYdLEoxIx
mp/wvpBd0je5DExSr1GhbHYG+c66HIPPFm6MdP8aLbjuNZdzZbzstfhmitSxZDafFz8ot+Jf89CQ
vKZ8wMDm3k8ZpCQNtMjcwkyNqNiUCMVum8YBv/1faS6dFpcAMuJoCHwn82fgULMjVPiNtovxqPRT
qlpgfCI+Go3FA5A1EdgRKgwiCgsomFvzzHewj6TFzn1VzaCCqsfr/1htln88SUW9jXGxhBHhYqeJ
WKRsb6zu03hq3R2SeV107Z5IubjWBTBlcr3rat0JU7w1HISkuQhgUB/nvb4Ax010kXIGmoervkF1
4pQMblLsS3x/K4l+7tsOCncV1GTtwSeEhb1Swrb952gg2hqvB3CGnWHwPvoiNG0GIx+kfKZzZrb5
2Yl+Q0WGYvtf4QTtXPkVi5RatZ+iKm1szDkU9qNz1A8SHxIXm5j1HVMcBpOm7qoQ+AbVGOI2QgP9
fNAXpEhjipm+yYE6lPMLdgJnnuFEyjm7gOxOSamPsrmuAzfnPgN2XjxWkXIwJk3RBWNmHqfo96Cb
NZR/HoUPsEJzHn8ggxV9vlC6/VY5wFRsvcCcH11iB4vxPMdbOL2JSfIkV5ywwhTrQP4qd5yie7wp
9BjGYCW4BOwPkj9nVN27GdgUPvEpqLXguWRonLLnaBdoHJKS1zJCGVhfQDovaB5FkAupZHjNsJNN
Csnkv7iKdwpktEuf5m2kZ9oder/LnOBehV7rSlLogiGDriCEtzO0M8Mm7HukGTnhZHEQ0exejAcl
AjKF1YGYqRv9nHLt9fUdRAFnM4ludDro21Izq94n/EyD9fIsWqv7OTTb9xaY6ch5v5G1ZtvABpvG
Z5JYaBx9zO3b96v59jTW6WCPlY9wVGme363rq+ahoQNNtXoNXmrVcJKFSKELy26uh68gh4AfKuwL
5KFRQfWMju9XEOJ/pdNlarBgIDdZO30iYxjAgAbkF8r9PvRrXid7WDWQtqy2TLVDpHHyl/0D1l8J
yu9YMgW2Tk5jWSiH3NozspqjCNQs8limfOY1CsjIIG6xfFEXt8nxd2DffMk8seyWRgdjbdf3lynx
fs7envX/MvHDiL0iAYcEuVve+/wCylk+nd1GRQoVeyItaYdxxvZDjwOuHHcukQx+cyiApfkBlwtn
mcn6X+IISwlnsYXkS0Xh8PzceZsDDNMVVSl0u170IvCiwFQ067BFPksUhgt+Jx6EIEIdFdc1SGBQ
fR78yq4XrLNeQYsPwBXgtPwuLpAQxCkah5wpm+xA5ojr6u+wkLiMcBv0RNPC/xORRgY6IVb5vAK7
i86NNpmjxjU/W7fkmCG6iWH9k9DPpub2yRgyZvga2W0d6k67nBaLS3QYl1/uH/ocU4jEnwcgJUKz
sNGOw4KjPzLOYN1hfne5Rk/aPJ4BsT3eSYXN76mYoBteFs0TUZ0jq5DBU5RrOToasXgyVdnCNZz4
euJ62GTPKtdBAX4UeceYZFbKhMjO2zOgq4a6Mhgcntcn5GeuIphGipNesaFPt8fC2mGg6Z1RqPKx
TyheWIJO1bZw6TGbIhI88LGzNScGz0CgbUusR8HAgcbFAOVNfRnsLolFxl7LLDijuzC1LJV1ScvE
z1nOEbhQtCvN4yehsstAUm2yKENmt0IMp55mxbVkUXjEQmuKA++5uynObRO+56dsdkfd//OvlPTc
ssiaOkl1i3Qy4DW67NAp82wTWbjD+c4WnehDZl8+D5cgBzD3UWcMv/qflzL7eej1vZ/c4jumRYt/
UxvzQoQHG7kbysif4gWj9Oxtw6RZeHERJRH32RntBblwTnMmHFFaWU3dcyIyIhpgRGsvzDcSYv5c
aH1eFIzMun5qfkw9AJc8hzyQhaJ7s2Bwyc9wR6zCiiwpeulupBZ5+hMJU33EoC7brbuyCOOOYKTF
hXuYTANOH0fsYQZC8umlX8AgpkcwBUUea6O1+kim6Vr+ymBFp6Z38hSVeRkNhay4HSeCwmkzM5H7
vwtkZO7DTdkF6xXgMtoWJSQDe6D0TqXEYjoU+q3nm7PzRVvvtFY15PQ5V646YAFg0cHYnUCcu7cV
kZmRgHGO4xVIQ7W6PxVIqfqm//N0CyaDAXqT16ldToZVbzEZEGv0YdFW9mioSh7EtsYzJ7Bux7Dn
1U53Mard4CZIiLNGgVPsip3qyYNdp0bAEIJQtdWJp0hhVZduMJUO5mMM7t/BCdfUGq6WeFmPtVnx
KhRPGiHIOH49yTV0LOgl8Nkqv9hf9E3iCqjYkWFjh1eBYmMJXcd/bQyqNQLS5KtPwEwCnTSfNndp
26YumWByw9Qrq2kBmwBG0ewjliUA5fukiieGACzDhAHro6HgVfh7Yqe88CcP3Cqz65Tb7uENxKjO
rh2vPeZwSXN1vj84YzskatMkUP6WHQbuKmiLn2B+/qUN9r3+22O6/H0DR/q5lPLp2qWxIFkfKMOZ
9IS6G1mYlM/hWoZg/Bk41DFQIAhwxRrTkh9ng14nVkLwjPu0F17+JIMke/LUceW0kh7wVhBRIDf1
huOnF1wwrXLiKLn25yVbBPz4ljGfmPuJR/hVjhl247MtuFqzi9XKht7so52X/ef3pSyn0MvbFLGX
Er4KwgKQUoYjvrgd7z0OUxjN4AWAFZdGrLuJF7B+Y07Q7PUBj4CShKc4vrpoFas6HnhUBYRiJz0a
O9UBUirZJSoI7rv8UeeCYEkLKjqY+MFHfwtrFpRjTROvw8qPHn/qTYjk0UAdSIw/6gWEzT9PsDJy
w1aXXWBmcZYZ4HFvmtH6TZ1lk6UpsB0M5xzR43vC8l5qa1kCv0X7VDlPzBhrx/14WfFTBQji+luu
1MJjE+1Rzi5tBlBBaKp85+pf723/HALfFW8pAomRLpSKvAWeCkYLdwuLqhmHQXzBnaD7EqCHwG+i
fhH8+b2TDkKkUFeWJU6fNa0KnEQYE4evUGGX480Pnc1GvpH/OwHpQyxwfw8YM8APb6mhcEJS5+bi
9BdqHvYQbypEHA2Z4btyTsP9pREXLgjStvEGW7Tn9YK8ONVqKDGOR507VBD7b1M1syrST47XT03S
mmqtQRmGWufhhOC3U1UZJF+ZGJmH5vOXiJkdwPK4Ipm4bTEua4EEjM3i7+2B5F7QXsmwVCvkhAhj
8mPjE8bXqHi4FlYadS8yxu5ZPAoJHJzsujTvntmazqaUSKEFVZw/TdY+szYb2FBeGlyNN6Ssb1eJ
1NJVXwXLu1VrT5KOZOuyKh7JIH+gSPckC+64f/eDELxr6pvzaU1sZogmQikL9yW+l3YqBrNNl4q2
tM8h7xC+7c9CHGw/b6ygUqmj+dd6jGxPDtUPcE/UhcIjcdo+yPPV2EHthoJlYW8FT9SrlxBuaGLE
Fn10j4kUVsb/HIFEWCp2H4chzUMVDWSm9ZUqs5GR8GaWXfVnHUgC5pBXSF+sXnges9Mpp0wFqaiC
g33VZLBPUwf644okNt0vPr5IpX8hKnUvUglInI9nFZoz8T3J/NaYwBVcNf6zt1AOxbyxUuJvRgOU
8KbQhjtzIOKUDHude1aR6WA1WyyK3RnOfzlg4O8byz68IgWDX6/eQXiW47pA5l4NbySvcHJh1tim
Ju1AWXxJbtUwzf9b1SYf2hvxPhSEC1/IYwyaudfTpzJNKAHnH5TBTREQXjLRXr96EAcY9UqMcqLy
6RefQEdJF4K5i+ycZ13RwFb68sCoNwVJDsMhS+bJW//APE8nV/r63ZUefEhY8mLoBzCTa6tCoeTf
mVaHo+uoqreY8bzxU4xEtOVOJQwZENeW25p9Z60Y+P9zfPZxZPbdcEKalChzGZsql6xgoz4sJfar
dcPZbqbafzMYKL9rQONppUrt6Pycy0UK459ieP7I/0FgpAsItihQtW7TaRln/7H6GLcQSUhkA2JV
UE6XeLv0wPh4ZNbmkJEYsVl8KQq1t9WRx9DDx1QqggGNW5nC1eFqWIYslpmmT5N7fFfLC7i3MR2I
5oGIli22UxVxLJJMv1QLMC/Nu0ikICUYtr3Kj680Wr7/UmkYHTme8KixXys0+UI0LjzqRvCybWYR
tCDsKuaYxFKjsNr1M3yg7Ljq/FDGD3jYjXnrUCy7LJM5vCWx3G+OXB3pcIkzfWaVk8k/yYt38zey
dDLIo+hSU/swe+N7igXViA5jQAwRH0fNZ+CmYnXaQxsY1e8kDi2PxBe8QNDnIp6rYBng2fZTyPGS
8myR1HAdgshCdSvIyo01XtNWtolY+cNrf6vt3Lnj7KysZ7YrNUTVWshysMyz21UMJo114KGGKfmU
XTdbbCV82BsXOKJPbTlBp094yKKic9Mld6qbOQ2jO4py+Zb8E+gVpH80mMxaCoSB1H/8JdwLkWta
kLaAVSxGZ2HHozA3mNzkEImOxUUg4m+OYv5DdoXC3lZB8Q8fxtFgLM3xD4TkEP9NWIp/hmmIETtX
222xrz4U44LMlZFxpy7Oo42QiLR9fYvoeOH4Iv4p10edpyLVeMRhd91m8v7kCzuzOOAJ5qnEco3Y
8rt3qmQ0txdCWdDyY3X9F19HZrO1Dkq36vbnliP55tnioI7EbM/PM4J4bbQELQdUMriZc/1+1rf5
pvQB7bsJquq3szWuOwMKSfWFIv0+q5rO1yLCKGUEeciPaqhhF5qk4JD7TgzX3Nt6LKHn66daf+Jz
aH9chXO07Qo51fLRYMgtXcFUPaRCYNkVOw4+qVhM6o8bgyVfp1sN9JEscF2RThsUlI6HeGp286U+
Jmqm4R0FZ68O7lhrDaC7Mq91b5Zbigyvc3VnGxXNMmPnzShYJRHge9pwUbhaiHvljq1BlsZQLkll
tV/FIjThG9mo65J4aUYgFJNMQfHHAQ2WFWyb1ALT0SSzVcoUUX8j4t7KebsB2+L3R3IlDqzbqIBI
HbD//mDDdtH5rRFeTutbmwxyXgAXycq/YpwsRY0Eh0EE1MCwI72WhQKllmTFHfdu6ZUS09mam9bW
uGvMo2rjZeeo+Ja/lbBtinBIu/bwBp3cO0BzosOc+7ye5LEQN5x1VNXQtaolZLIZWkm9nSdHvcR5
yVb5XxPBrkI+QVaQ7ullHYB3yFNmjdsSbWQPbRRPVEaRoY+AQnf6ud+AjA9edNYs+LTTRPspYqJQ
GhuoV7PPIRabQp5Zf45+wF4RbGECNPMSHl4iyiA1EvssHXs0sGtxEtTaT7O2B0EF5SGNk84NWQr7
ljbHaGIN1wfDPgu0NN7mlhR+nbq4Ha2EzSAelsY1KMGHdG7TXqCF4VDkwEKKfzwJr0hRR+34sfUD
GwE1cfUJV1yAd2Ya/URi2HYBZL2b6BVTbBHs/73931cOtLxMV15vfuCv1BqhDsqKbFazDZU9oZQl
GgRgVYeW7u1Zayh78PpmHciLrAslf+fBwsLyWo3Aa4Vzwit10wAvff7tTCyGY+sPvZCjC4oLYe9V
gBDmVFlQFY7d3WwJqnZsRIpL3MStGb2wjoOAhUyimNEkIJm7HqRSnycprjrtUOMpZ8ZxQUB0yGEc
vGbbq7j9LZdSXcCliObdq6QcLD6LwtoZZUUKh8uPotvHAocB4wbARI5eHGb0m82wqIttKUxfdJPZ
B520x1AGDvxiU8DrjC7fU3bx4UWwSEj0zRs0kpC3qgc0yJzgTqlnEPAU+5nbizn52ZsVcTCyYzM+
gjeMx7CkLt5Wr+tl0whX9QLi7CbkVb4zQ6PuRBejnIFZYZ5WzNEf60neHzK7/7Yp3jONmtoy8fHO
lC+/RcCvAWeoEj73LkCIOK1bAK7neAijcrsg3SwQ01Xqhqu3fKO75TuUlefsB4niImHU8+5Nd/Vo
OzWwbUdd2B4lEqJHo6AEqtVRwAGQhGqE0Kys3R4KXwORV76wGb7AmSU2r2Yldr9rCiKyetGs2SfH
Wu+bt6A1AOM4TseKGMVRx9/r695iiZTpl29q+NtaG1kBSuOoTDmGpMOFF7T13pTiMhcfqSUQo6oP
YCACon3DvIAVSYv5Sq2ZpMpISbHWcadrAqLzozcxBtO3ENy5GwsSt0fUSWD9DAcPdnUI5B97MJ4I
DvrwVkKSw6DQLrRVoy1/plcl/hZXZGGHgZPzhFZXTCV5VxEIu7Q5/BBM2M+CwXQNH/Qe2oyOxJT+
OZfQ7rQxWp2aVY6LqVagCF6mldbkQQP9SLIzZBZ1DlmE7vEgdIzx769UKOyQ51+P2g4EoKaDOTZv
jcjP1bxZH/m3gl15baNWeEVB0UjpgMUdL6cuthEa10/sjm14qbdEsChNv6R4gItZEAMv3gMAvuGm
tkDV+Dgtr4S3/9RUTSg1Uv4jLzlyqNtc82mNp2rQRRcteGK/9v8disS8V7Q80dPKCsv6fWzR9ekJ
bvcTqnZ46o7yMqxcHvt/UtG2EinkPyyWOWpzP80R/8CltuPygpROwQT32yq8k0bIA4VW2ucuymIK
MSj2nIbfO2ehmENVvbZ42q5IE9oTW5/hX2du0ZZU8kJSl6QVIkqL66Mo9mF1JtkUpMb6HLLAou8l
nl6aDgvDE7njoQSaQA6y5FVSYEwedGIjyuWNFxd6jKvVXEaX027bjNClsXOpINdB+31C1znQHmkv
Z/TIsdiljxiYbt6GJBh+eq8I3otcyU/CvUrW7/w2HRQrRQu5cVb2r+Y7qecTBDMjouyBthElFfpf
9SA18yqYc5sUGq7IflDMIc/4HjZX7I6z1K8VUHVjWGtLjUHwnyLmXaadCLoccKZyjMG4brHfmgax
hGWkgyCYEMkXWwNKw9pzjnqJkJ2r2JrtOTc2T9B+rYuSLrgORgUnuNDDp6zPVObjgg4P4gOiGlHN
H1LaxGec8Es2+eCJ1M7X/54Dxjrf5Aeh+86954oluqSDuuC8PKVxqVDvXT05geVbDq2AovQ5tU3d
D0jlfTI+jM2F497+9TO3rJyjkA+KA0nz6ALhSZYUItZCFJLOkY0Pgi8WDBJFF7szhGD9Usfw36Hp
7vOlYEeO+xK6AKpw6wfsrlxDPTfiGPhUokGH+Qb7ecW8GriYSG7pUrOOjk+HDM+ElPg6ZXpawvwy
QElsyIPZpZmC6RB+30tmyUdp0t4m8JAoCdqscZxoHRw9hg/CKtuFt2MSXFavZ5r97D5bV/TRbsaj
1bBjXHIzng0F7xaNJOz6QeRFOVZUoZNMwNQzDPZtOrChXL1Ct+TLUCa9+17RpsFtQQhYeRCbKVWd
mhLBdNF6B9DZvzFRi9HzO7NHNGt+5gzzC5ByXEnBXf5sBww7DNeI3/z6+mhULuLx8039K62iglEG
Yj4LwIFPvp8CEv9nqiepo1nw10yNZ+Z4txSMRHwyxHNyY3q6DAY4bMHVI9HDu66QONdxKMpHmvdj
dSv+EIQbK2qWVCNItMulnq920K+4uj/CRBucgtMei8ncgYNo2ybXTWxZv9aQGrpwFVjuHHWIzZUD
HDKsXNtoggF4oPRp/KRg/RfLKXoqkEMtRaIclXs/sZeGAjRXqDznHNeYjDOFbKTwgXPPuzzIdY6C
JEa4GRQ4fpsobKLy1/v7SJDGNYNr7xJPmaxR6YWAu38SvIy950j9bHXFYTEUWO7octF40AIHI/JF
P+Dh/k5fN1dX3ootzKNzdKbqAww+aDGD3bXLZ1XfeN9FHdWBL91DQUQLLXwq/mqBxvEksCGFKfPr
UK04JXG+ZRxcbq/5hJKhKUQxA+eyq9tGqoHq5KUe3RL71ds0DRYxys7eOuQll9NrHzZx9d2sVAF+
pejjI16zFmMzNyC4h771UWCY5P+QqugwV64KdIV4Ckqb3Rd9UAOkqM+UT/T+gmhGYGMO/Khu/9ls
57EHd4HPf5Lq6wc9ktke7PYlYOOWv/skMXCO7hTuMGXn0/OyQPzZ0+/L6WMBXJ+cTfXkdwcrdXX8
RyT18ceTrjcyBo3zMX+156iI0E5U0N0iiuNMZNxDA3ylhPknhHzxsX6yf7BFNm/DVhwWFY/QEVH8
tiNUY5ztF7xaXiK++gSs/dC7yXX/br1K9TgIOuGSFp0ne4Wlj1bUu08995T0XTBqHtQl1pkq5Glo
wXIJPiCixbVqkollJEw2wuIbil655cNUpMSxA7P0h+b0bKrrZyzfEyYSm8FYEND5xqfmKecSn6gZ
1uCLXjIBzTl9lFyyA0tFuNbEFfraN0c4yl2awgsc1HdfVwB6wR44JunJI42cusC3CWBanvuGFW/m
/VcW9MUQBq56cVwyzymuF1t20+bioLz36nIQT0vKN7tYTEMkZo360zlB6tzGe/1yMmgb8y4ScP9d
0xplKNq0DBFAHndb2YQKGOk8WyOeuPeeqICCB1Mp50LnIoFAYLCGSds58Z2/h6TYCkMHZOyxccqw
KH2R81/LZ67yyM5DezF1vMqmTMOtwZXLBrEY2YWEs5Tpf6y66VspTiA0t0rXY6T63ugy7VAV+phb
VC4XsxbvsKkAg4NTDN8eSIAx9GpCQn8nKclNtrg02+0RhyVwPBQzyt5vxZNiv7vw9LeXrAJ0NJRx
/+mDz7XOryILOSDgUHE7DnPUnH7MjCIMZ2Jnph+9k6ul4bth9HuyLDtoJY+Me8RQXd4WZDK7AHnw
jM9aGv6l4y1pGsnp2drlhvrARqUP9p3+HZvEhaoQK1hDSoYBEvDKjdWCj9q2b1B3AuPf2X7H8hYv
kng3wseHaYQcwbNqeenTdiKCONvktLO+DMsJbdQdP5NdvWqLxImBAB1wSz9wWgUsJROCjrnQ8WoV
tWXMoFBp6+70mwQ3icqZCarOsJMd9waQiXrKd7bsK1jn3vLlSxP5eu7kubYD+5V49WJrUh3pLB0b
aEPsbl+aYhdDPyCaGsdB24lQaC1pXbmLeD+HNG+pK0xN7/5w9SLxwPBuxYkLCUvIy7xBnGRWkFRw
h6Loc42yqRUCqC9HErlsojXuRb0ElwDUw2DQC4rrc+RrGVrmzC1LWBnHGy4kgdqwYEJVJBed4QLf
Er3x2c6NFQTAUcdJTDi3ud8m20FEBm3TwhXRHbI8DMXk5e5VxPRBa2vRPlIMtUFaB+MXBft5qjv6
9WtyMnXzbMI82hmOZpteiiIHEN1pQGLGJG98dEWbiRx9rx8PjkrlKE16/NJqP6t8A7SPS2NoeUZn
W7+pMcl7JZBeb83kA7q99E5uZIQPd3OpDSA0Jpa6B9jTWr8VE6EUTxIQCyePXkM5fR0JZMkTU6rK
HBGw5uI0G3qjBRV6dM5sLpfrTgTATdmJHFsWYhcaOcOht1VC2BCUOxVgcPk8xWLRwW5pAOpnaLjT
SA6gNbayj06l3EbwpVdXIyj/oHgz8tDPVrLsoSP0E513eCdVjEaWFqmiPrQwaZEt71qcNQu5X4ts
6IycR800YfwivxwH4VEKLlJxuw2moj5mV3uSjHJpl+z0Q7k+7aPaFINTp1/Y0pwijKveJrwxcl+P
Sp5B0dAi0qS12LWS5jI+Ek66l0aOzSeLLuSaXEXam5SiWS8hM/GkUwL8W4q3lZ9rFOA7s7AjJvwB
6wjFzPBu4jRaYRjutYHCRApagnF7g0aIWUt8YKvmNZDoBBd0oyo3ND4+g9bn5TRn+E1tOiv73Trs
AIkcNBx/QKiLGLC00/upG58cbPqritgHnYwDH8sTvVQ8uDJ4YxFF12ixq1qkexYg1w7+B3B9hW6o
f/6zZL4OVOcFydSm9xJ4mNQu7JdOusm9/UZD1cdVNuIE6sw6x26i9xjjFfH4laxgR2h4Y0DSfFHn
QwivAHsbPf2mUmw7x8YHwznpP3UQ2xVmYvx0xZUJec4FSRW2SExCg7W3oZsus5zzdbMO5844mIEJ
Otngig4BskeT8CrXsZ4iULc0Mdb1CmgYtmfZZ2IFlJNHXYRn7w27fbDcJybPS97Ia7S0H8o/jjvv
dvXQgyiejLkZLBcYCZe1Ph9fArm1yJOWWaYZkt3eXR0DmYSfyvxVIOcBLli6kxck04wmSA+ZEWKa
Ib6kp0x3h6j8p60Lfj3H2xhdItGtgRk9Mh58VbN4EeVYCUfIHZXnTYwypLaGqgbTFA4OIqnRpRVe
TKFUCOJt4oqACVEwYnPqkd47KQeUQd1zBj5fvVFC6U9vVMsxo3DU0RFE5goJOpXVsSp3v6L2HT1t
GHd06e4vs/R8bn7L1NE1ecFhHosgLBb9B8Y0nC/ndgh7b97tqDzp9LHc2+zNkw1hfwyiBxw412Pr
HZABWzbz7ysgsNg/IXC9iWF5KOYx/YVnhCOEzdXVM7g2j341lyQt2eNy4trIM8XSLxE0lga5pOva
yo19wydWCTXyD6Cbkr9PzC/AZpr0WECcVYTzgB26nW5hHBk8rBugf81IY+4fLULmUFCxnhTKlPjB
ujNkLdkXWHA/p7mZwnYqYZO62/sRzX1/FVw80Pb1B9AnjB9M/myWoKFOjaNrgd+kbZveQirP1SBo
68LmOSqMAW5+uxpeRdUm6B9nPa8uT4DCvTh3F059BwaQnl1TAra4wCZlFOEr2fiXqAIusaMFCn7j
cE/8Hlo+FW9DlXN1NxZOtNVXLOU3a/6lSRGLffCJoucCiEs8ppTjZI2sMYtSXShzKero6WqIykrj
xlI9HKq1zSnU29lrAmYeRN1du7gxBv410Phr6Igyjw2DIU4LDBO+ZbmiRsOiMhzfQ76Cf44n8bwG
aRHfl2mM6wmfddAYJrhwEWtLRBJh8axtOUC7/Y1sIEn+g4iegK0bsnm9JiKFRn6QsGtcCJvv6s3a
MvzJO9IamQyHUA44pNMeB4bF3N7QXGOYoZ1/MWmA2F49Lo0DmbPF5jfzNGWWw6btC+HzZz4iZ3Gr
hBvK1vQM8QrhNibThlZLzoYVAWw5+g1UiYSUpbNnU0T4y+fxFSN1YcWEr3MzADkIo0mgdsiLIBCB
sWcFZRUACcCOyqhAibo/+zL9VKgpyMgQwrb4jXZ7F/fkTmBaTc4fbTEh8pB3kRZJRwbKoqXSWnsl
WJSGI1VWeTW1eR/95oG4Bh2c00/1/L2ndm+j6aAwU5M00TmPT8hKRQkOGtnI+izzI80Bar8TPWmf
Cgu1qecffki3namyw/WPEd24sBd4QMo1+glvlf+TPB2UsPdtQiiZ0qgGIZR7go870rD6pjAc4Kvx
yYtLushF6aZtqjTHtifyAjXrb90FjQF33BTkxhNU7+TptWHlvWMxVaNCuJ/x2NcFtQGnqUeUjRKj
H0OzpczaqOJp4Z3bF5A8SLwC1Jgmxa+9VYrJYGgh8nB6R1R1blVuJAzPnX0LafS+R0LWN2aInzEM
jTefXvaSfEzfrnlqU2PlktXRuhlvNpwHhSzq0fXeTCuFLkKyVSdr7Co8iAWchxZx+hgYmBfyLBr+
o7TYm+U3QyeY98FrkI+FYcRYdJNu2xrs3g9Eyp/BKDQxC4J//GeS/4OXSMoZHiJ6pY0yxlX0nxiX
oQMYomfWvlU3AT6FQDbnLPcqIYRqwUsHsYQ56eCfBaz8Oph5RvO2w6bSH0ShJ3po/6ILWXuJON0z
nN84JR1onDbKJAAos50qqzJ7fQqmep/jK1p/EHxIrDVszBsuCwwtirQQrphdWYvNFAJecaOHaJai
YpBa3D3vIaKM4MYVBQFIgivegUvJj5uvcA64IvFVdmHbQZXh9Ozvwm3apsSuQLcdsFuHCt2Jx2Dz
Z1EwMdDL8A1QnuFWJ97PvrrPsUNL/LTU68T8xI50dpF/OYvox88k58IGrEf+P9znHSyoG67VQT5/
VfnAZF0j5Gc3MhWbW9qkD83GyyMyrlJLl36KbIpEcYNO09SxkPxsp49KtmlTRQpofcmtq9cALZAI
L5WIz92tuDT1NgydHkDc/mAdIMUmaNgVphutVGtIqFG5Ck2Wo4MNz+mNTQFGjjYK0Ff6gJB1Hr0e
uB4rS7zZ2fKn7AZXIkPamIGuFXnBtHaahfg+JyfW9CARskMwCFxbDRuUGVhaTOdUzaAZ8jE5DcLo
QtxMJeOEnlPU1KzJ37ZRcVAMT3YC+dDt7FcS7P0Y75XPoqCqW9DivBt4WBKbGkPikiU2IxqEoom0
Q+iShqrXnC/hJlQ5TA+RHi8prQN+a+iGHDrw5ivsUH/8qSzR3LJ62Z10KHjAbQnsXYmQrn6tUbuJ
8P+PcJgDhQJaXp3cR0u0j5S17x88YCQTqEa11ZeceY+HcsKby46Ymw1jNzB84pPHoGv391PZWE7s
m6uRQrFDtanNUowflI3D4akpOKEuT+q31OFEVibjDTsvYvTDR8HovIuov3N1xVDxmc8Cwy6IiNh6
7xrzKEPvLAEL/eHdbiBpDqpBiSLdYErlf7TdzUsRhM+zZRb2ozavW3Ml3MLgJ9XDx5DHcNfKQvvt
im0FHOhTgJuPU++JI09PjPRNHWJ3u4v/YXESMFUMECDkYAuEYqb3vk+TDUzzeUL1WV4g4vbYdSlE
KeZqG30aouomMSP+bb2w1O7Lyk/h6tG0CXm/QcvrXZXtBJEiL3fCO1iBe2vuW2Q5l5fephUVR6Ui
CmFGmx7rjURUIZx1Lpp1TYYRKAdfqVPZrNkbaoqD3/KNnagQ6gLuAfSJ5yNSgBHZLkhHt8P9R2Vg
mLvxJtjx9FWlLPQOKYrGH8Jzimd/CSZ4LRHBNc18R4xfNsmoFCr8sFTl5ECVexK/JoAmLOnTo4KC
plkMDpXtLnrpnxWGU5YlhgGNGJboHD/7kNoEYaunWxYHrFjoYtwPIdt9QeGFGf6qRRNZxacxZFmF
E3W/F3IbJn1nMa6dL8mBDuG7zExECmrwjVKR9hCGNeOVpQIeqj7sDm0SWwAS9aXwlKLq/1kmaeuI
PmShdX2r0c7FX67c3xSXQ4n1oHmyZMU3rYOb1KPk4PpYZVj1bENNlPDKnGLdLhxL3zM/6zOtxY6E
IxAcmvf7+k8a1PA5MeatrVQ8WiYTOeuPwRCfDSuMTHYEjek11nDusUnv6sSqi6uHuFkPBqT4OZl/
25C8z94jAm0pus4iWCRDvnwZ39QzQXWv/AdTts9jMht9WnR/4gfoJzXYk/xYzMpZM2N/CP9W+S7y
D5RtfQUC52tELgbjGWQc/d8gKermIBHo2hs2TCh/48gwkqmJo2DA+sEoIUSVjJ+4rFmGfsBnuw3+
nyht1rkCXBufsBFIK20mRcihK2lY98z7zhyKSw/IvRMujyJDka9F74s5vvP3uEdhJW9yionfGhoe
f/dhl+4krk/mVRT30RpwJKTGpg+otQPIU/vFQ4BfsOvZPPt9Z0ykCMzcXzuYC3XaDtf39Svh8J6i
A9EOfLyUEXAk7nMslXgPZLWWS/cnn58o4/adA6Y4Q0FbKsCu4B16JZ9Q9BPFW/pBaMj94Hg5gulW
ECLQxg68ptD+lgx0XYsHMC0+zO0UqnjcyqK4OKX7C7Y234vfkbqY89ETYNtMsTnLFco6HHDi3s1p
Ip5u/VVqtq/isbFtxBM+ViNVDNER2vwzx9l9YyBSW+LQVFsTg4tELbAQHr72iNvj1XYc+51fCLeS
ZuSHbxalUTtT+uyYGL/JZYL/KKKpANjDtKMSb6LWPLqANMF7uNhp3FdJIP3mglqKc05L8wmeziuY
QZ326z9wTkBYwE3zt8UtQ1lGcIslphubehuPMAj1phs7GgHaiQ9dRqb0Oz9EzH+P/9AXDgtnfxab
1GT8qYlcXnhJJnse1T50h4OKv/Frnif4o1y9AVXnsbCbSf2yyvzyopcqakMxJ52UaWH4KyjhnNuw
ce2BLYRhcUm5VxQ4UUTkcUHS7o51D/vlB3xm9QpnpMxZflWzp0HiOR8tF2QXAxdRJtOO+b5vVXU4
wffcU1UCtL8VVxg0W7Q2Lg8orFL/VYO2fO1u3Wf7xPHSPnL1qYPNguAknXY6O5f5jw+vxIyuulqh
FYIEuLZ78yR7YV0SP2VJoyrAinbhpvy45iKXfDacJgQsnvYRUv3ixOaTNA5ssHulnh2ViJb6v8CA
FQMlGM8nXgonQ36AnvoMRlpUiEC7YD889LmOffL9bN1XOi1hHzjW82Q8ECDt1aRZ+O0xhfSqeJII
/xcDafYQanV8+xD9frCFEWeujaQ+9UNLh9Uu1jYsmISk7sczwvTLh268gjPMtHi6rvVO2LUvu1V6
QHUihHzNElOHdHj/S6/4lsp91E1uhO9IkD4MPbGxjnE0GdNnX+dE8LKRUlY4/R+bc82otiPiS3J8
A42GlbuqEp1Y3a+z9asgCXQO3bb2kIRtkWQenW0XQwBdqO0YxLNRdBmokn82NlKsO9o0X0ri/+mj
dshN5MCzDo/tI/U1JfiPuReO4k7Fn1AlJonctMRLYodEUPVBg9rn1mqAbIZnXiVct6L1MiE1KVfr
b6+dIqzXSbuWoaeQWet9PRVzbw3oGPRZ7oJu6i8HnvSOkCrQxaVENtwh6GV/AZvNwGo/WA7LR0qI
tmYw+dwOQ608SOblc3BNxGaVN/t393rZAwaNf+OK+uNOsjDF57553mZ6/RIXJsPtL7O2+vSh+z0d
aqPbwnHlp+ycs1DbJ7dFEN9ueHWbXoYX7faURZg4W8EHHyC+RyJAjH2/JnFAzPhPWPNsAHt+AyHU
8HPrlIRxbvqEheKSc3EjedkQVhhu0Kz0jH0Bu3/QBK0abn2vB/KbpNQXC6Ja/RGd16YJSOiOFpn9
DYDegyw76kK24dmesDpN0h8BdK6e8KcKZ4L/LIzGDD2j6EJh1lRQHf6GVVGPxGrdAzLTyB2LcCVB
I478qOqzP+gig9+/SP7FnsWpYKqufZqbiFUiHLrE6caTcQQiCGHeWEzF38Qqikf4BdEbiBRkB3K+
ddRJDuGdGHPH0X9C6bGSym5kk5c0jue9GWBi49dna3Ipty3gP7K0a9QKlJDJor9kO29MTw/ZAun3
1FfOyTlJ6EvpenHZcOWMy+jFawv71vAtZtOPN0MCTVDkmCOB7TtIy0OjAC+9772iP3KfBMxbs2/8
oHtJttLzNHfIc6Q1Mk7wzVqSpaV4nLawjDaHdZqmWj5BJ1h6c5ADoMRKxmMHZs05kACMiuaq1ACR
sIVG1MKy9QLG9qDbZ6QJwNQMvMOf9kInzMhC1ae5ZDtdTObDK3H/Zubc3bAigAJoKaOR2daszGzp
hpgjf6O4Gs/Hf66w/BT/glh0cYiA3HsGWzA4rLn6MjpNWFHV7t+gC7HzLd8E/Kpu2nJsG4Mz+HAz
2YwYNkfepykJ4m5xQPZnjqxUU5qJSGEcYbijIjGVEsQu7DPbnRn5UNx19QdMQSei/kuibXTMRmZc
h2N6eKLw4OoE0ZLyFxoFOxJuA3e34xvdZrlUP80AnBqmCsv3yOlwamq+IMOTFf0SFqIwdf5Fgbfl
7E+GmlEA1Yx/9zhPHXHwlokyTTgVEJLWwVC7NsypXC9Q/gh6qPrTJEuc4e/7bWSgBjt8Vfk/NRF1
XQAmJ05UiLxnmzoxl81U6MvjaI1uaoRbGMQlUDLRLRcD8zSRPEfHKFJA0/PiLyJONeR8p8adBHSH
kZUCiRlcBmVatWNI2yDG1YGibcNBGJQXbDymI65gf4MqIwH6ILw+k0leuc3luTeU9mobFPzXqNuF
VkIN7yA+9/unhdsgzfMBKH1cN/wvI/0NXrqQFRv8yApbRAco1Dezfssq39j+xwv+X5f0OMzgRON1
iGrBJVfLwIaxC/fT7eUD6/Sk/UN6zvuUsqktvS/dDPGRLJ89I+/sS1VKzFqEyCtZnSLwyoUmH4nc
PqeFCyNbfZxpIy1zhn3NwLJI+noNDEtMDBdheB8o3fG1O4PWyhmny6/KCGkJ2IO1Kr75INKRWJQ7
xxFZfWuUiev9u3N87Iq9DajqBqtexgp1E7WHPYaaSOKQ8Us1hi4DNffi7vsZEwYm6ObKV9IcYSCT
bmDvibUhCv8QASq4LUW8Di25+Gl90ITtahcLtNF/T21bOoKkISbDFrUl3tRSF8xqcqHBPjJiAAC+
Cw2viIFQlOwZ+l06H465UwP3P5SEJj2LoRdTaTW5sEmL9ihUH8uS5s3aJx8BJDiKNBSUpbnzJqev
JylhhbIvoJGpyHFwdUlW+Rx8d+sFxryIULT3UDUXvB1NmIvbdnFudWr99nTx8APjGNnDyYB1d0t6
23uboKSO0/UqdumQLQ7mRV7dBL4Ye6fEiC7cVMGRsXWO1tToig+6FSmo7OdKQa/X8wudiiMlAQlR
X8WGp/2Uca+ZqgFKMmXeBHKGkF0aLvgF3aaOLMZ4w3FqhcWG/E6IhfyQTn3XfR09P3PGzI/IKOBf
KWHDJoV4Cm612zz9PH4u19xG6DH7vn/6287oMMGIMEC/UKgoVY98w+ttH8PbP2qZjsJW0I/5xzv/
Opg7f7Ic+gF7qdTvWFkIuL19nceSjPTCRuBZlo60NmOI+BJP108zk6V7il9K+07VKtjKr+zSKImy
TA64rZy+DinJmG95EGprh8S+7fhjqA8JOYOdVsWHwmPvoKCW+fAMm1Ac4Nm0GnZXwZvXhCuKx7C2
u/EhRdJdcyceziB5tSr5SKqKwaC8Tql/ObYSwFz4hyGQda3l1YnM+fkFtJ/DLmgUHi53e22OE3i4
IiW/Eax7jVhBe8MLPTgEzeUB09J/ObNUahUboq8ZyNSgfGgj0YpdfwtOkeAr5jHsy/rGnqQZt0B7
zRx7IUrWR/t/AHQmJnhDEP8j0PrNWsnjl3oVlzeAGD4yP6OMUZdd5K3SJDD8AGBmuZmkjJyeil74
R8uPZwrFuVH0SpFW+DfQwMIWEOnmsebegVi4V01dsmST0siiEaExZdS/q+GPztRPFJaIncL7ISJQ
ymBppcy864/etHCcQIsgQiO6mI1UXYdi0Yqqa3Q1NM7xzlBfBtpBa+idi8bgLcRPeCB9tuyiTvh9
0lOg1uUwMP0lNHqs7hpxQWudbqGIIrh08QxEt8wLzis9z42rtLX3utxYKonPTmlDrE4VoiWjIk0m
LFyrXhHPkaEXCv9CJNDXEfN4qdyzGi/y9TdLNbfDdKZv76X0CUaKlylyb1F0bstWq+3b4V06pB25
RJh+Z+NHp7JSGksrvXvCRaxves1M3r+cPbYBIBOCE+HFgTIv83eOmTL9SHGjZDou9k+24bKcdnxM
1pg1fzeNDxzmgmw5+Wnbhl1cLxNmO42lymHlrqwM+BtsDhSq2nqMA5ohL1hgPo6C0FaS99YQdIEv
QbFlDNpohZS0xBv4c/6zMTNOiLPzIvN5SY9pnbzAdm2frEf+mRyvBCmoDe9pv4uEozgskn0+y896
5xRirBz56yWp0Uf215YpA3Q7DJvQVRB4v+KVLMw3ogRgbZI//sfG6csOUabiEP/4s6jfRPtuTLm0
TldSgtCEK3IPyI9iUz/oMJV2peI2gS8WNe5CKANLSap4qYckLa1aMW9QRCIzLEX1n2nUjENHNdOH
j7NGfTCbofski1+8LmcyfLJxCo9mCQhxNDUchQheCdfnKahhVWOKWV9JAIfEDxbrfp36c3ELxtK9
/nYkfhXjVcrD5tVwINRir8oqS0A7A21XwVqGJnWl7RRM6tXtHaa4SvmUcouFcjZJxl8lHtOM66sa
IhPKCgI0jQRkK9B8UacVh+NNBAQqTtcGLzAsol+a/vN8hMHJMsKhR8oiRHPEqG3YX2/oc8i2Qlom
m7SZbHSJ0/EziInDiZHg0QazSr0iFv0QU8VDVg2JTkP+WoC6tBZT6mvEz5DabzN4+9NSrjQjy+fg
bJV7ZQFRFuKKC22e04G/oc8Dd5ne8eknIEqx/5lw0SVPBaHjdBfexoxvuu8cNQRQBrZJrctJiJmW
Qmyhq+hoWNyN49jEqRxvP9KPPF1qAT2nWeTKRdn8bnHvM38EnKAMHdoCSNVZPaspMR6qPECBSasv
Hx8dW/lnQdjo8J+825yZRqtVLYjTko9JcRdsC+pWh0KXaAmuvMMgNrp74YFaupM+ES2jmIto7tYT
nbq7Tir+sroYrsVUrkhO30VumGmASRWosB4Cp/KCGoINvAvM/uI7pPZTKFnMHd1hODpVoUlDPptt
nsyRq1ml5nPZw8et1JfF3d0W2w0fLY/S5gQX8rd0AZvP6ok3eHhCQmsnFAoupsbYI89oBVB4vP/p
Pw99uJe3JADqibKczRU6MXtCzqqbq53lO37Ob3NXoD3zb2qwfa4nHoBbkLYtz7aKwoHYIWmbadFa
vfTmjb2Qw6E2JvMvpuGaqToG7+Mq/46LlRwK+tKwIjNyNt/nUUG9h6f9Eq4dfq8zYd0LG3Gc+/wo
S0hh2xJsN0kW/dsuQxUQ9IDOWSSXSxZk8CeFECcFMuDbGb+cVHysbg71RiogjPGelK5uh5IwPAQb
VfSnLn2lDTbZC6TLqlSXL9xlvEd+68wx73ctWUPFsdpL8FlXzIgQgpj3TqOGFHvE2D3K3vo7OeLy
ma7ThnPEV/rbSMVOakPEqnCo6Vt8VQpvShA+SoAi2v6TnrQhHKfwyWvBONDMjIhxHdyIfLoFg3kc
msLU/VbpdeJH8Oaln8V2MDAUZibN8Xi5Kx/iTnxhsKE5eQM559sWfUqydFHZ8xo0zpdQt8eSfQMH
osIr2R10T7A43pWS64JTbkSZlcqCy6qjMzw20MgfXkXR+ZQNevXC34eoTAkaXRs+sR0kupSdajId
+iVtbbX/kBE4qr37HJTaA5Z46GBMoesK9HVd+eFG6eFxvVF3MMdjgkNpG6G5AWhVAX62Z+Wjvxq8
kDalyi38ZbeZaSOc4l5mrQDlsXdS8c49CfzEgyx20phoghFVeKnucjE+mrjrAcxk6JTI6LhVlgQs
Z4vr2brx8aocbHexSAP4Iflz0JD5ZzhYVH7Pqq5KsVeHLN+NTnpyxdgy/2Ie/+2FKmPpVFNCqqt4
OFlloAANGJWTbjirkXlOXtsjfAtQEuMpAykGGUfcqR4xDQKjIDg1WLG5ykSxkDM1i4HxeOkHHY+t
gXEDpBaUJOSg/WdBUIYQWiysiTHl1iuuViKdwphHyPD8NRBhFFf4pzpYvRzyF1AThKZphbKQHXio
4ksf/VX1RNLAov0WVD0HtcWco9/LqWNk6XSBMw7ih9A7P6e1Zx0K86V+Swbat2wnH7K7A7apLaiJ
4eseGn/9C2ZX5E+inxgMUCXtSC6Zc1MX4b5sPejzLMSW0P49WalK1+1lr0KPqile715CSKcL7fTu
QPXlLTMlAFftMVa9od3GkUb8RU+ycxPhho9W4vbUbaFy8kCC7zBNdQQbade4i7MgSe9auPU1Pyg9
kpYwehZeIBpMaRV3yrSOpCu+u/9cGDbUmrf5euchWHmt49/HkwBD70Fz7iDTE4l2VieYtrQaGWQi
ljmU0jNuJGw0ZFXq8reJObyzvoMBGzZczYRM4t8u0fOrpuzuWfz6yDruMm+aYPMLIL979HdHv/D1
fIh10sFEDNlqg1B2JbM3pkU9z3ZxOTt7BUwpAvCC5HO83zL8pWWHArFMRcxavhSOM54ZBog0ilgt
EeBlj22JJxrwJPo6L3C5v2sQ+VlU23GVQN56+9ZhqGFnTK6xTJxzKnEH2YQZJP6Ipd0BgPQvgX2D
91HTyIXKMj1W3KqfRyrzDKOmL6AvX6//Xjo2CH71eNyaFUD1VoSyrzLi+FTdH1HHb9IXjEjRSU0X
XXIKPY3LS4++TVKswFFSop38PzxHaANLipVd9OxHcenCZRw5lRzFgNKaT5GsaDJUZqaaBmbtZN7Z
TS3vNdE5+e8g2zReyBNK7V3AouAcI1cK6enGS5eZsocMn1N8yIZh1qixxIOtBDVDN9+UzGZlkwyp
f7JubVY4ttmlpOISgJcZbShYmkwRe30cUlybx1+Pt6wc0CXtR35Lsn2SJazA9m15mPSuPGlx+lht
9G2S8CArJnUl+3JvXqZ5RHAUa1t91KQRfzsAwPhtfY8qoNmcIqG+Yy4mnmo0P/YHodlY6XNoT/iD
CnFeaJsZ0JkOcs7u/ZmUPR+v/Dal0qW/l2oKtw6yGWb6lWyrIcKej7gj2hBpEgQ2QHY8ZkrHs5r2
RBFAUEBDK4ISpS1RJhCfmwSZPIFCV18cD3YEtUEI7U+Jc1LN3DBzKg6X3vgakrUg869aUtQiYP22
VsgEhb63bDoIEvQBaYGDP8X37HNeoUvN5qS6s0l9x6TeHMpqF5gNzd2rj4fvzRzNRBF3TdWkH6LR
t5pHay61QUMTxZybotwuceDwsIivwzQmnFBvWuV3ZxXMfwKtXLkVXFoeKepKUzC/lAE5429hcenn
gjTa6r1Po000ORO8VoGB0r1Ao3BlGwWIUmi2GcV1CHajdfdhRlNCMnhfuGecao+UT70Sf4sheAti
DXAzdeZmq4FwJ76CbDne9boTUqVwqBQzaRMUGH7WsrVh2lGElIP8r4AVr8h7zlZ1lhMssPP6PtK2
QGyI2pU/Xsm9dVTgz8t6EOy1BfBYe8BMEEk9/V+ITX8Ul4cWQkBuL86VDSR881z20eQTLLe88Ciw
MYg5BeM4yjEJgftluEfzKVO7WRlue7SBm28YMT6jqTJyuvpQG/ih8M6SLNyMkPfIFxe1p/OPmQmF
VObEo6M4RwF+9R21QeH9yT05BKjSdTkaEPqyjBL1Tby0sG/4Wsz9H2M5g929Y3Uc3l0auFxi/vjY
znNDbc9ZhoeAqPj0UZ03TX/cgGwazgOEQB6ApLMzIl6bAFrjovsw5VOvxABmSmviOLUr5+Qd1Mpm
gRSue8hvPwpbQdlaKvUUWAvbbcu8N733U2QkJldI73TX///Rhsu5hFH+ygO6Y4ke9uGkJB/ZRLXW
wPlDf2Oj7XAAoTeNmrCIUbCovaiiHQM4nFh/FaiYF+GsiYhp1UUAV5WDwzHsdFW+/YyJ3Vf+583Y
Fw2jqIfvOu25EkB96+l7ZFJNjlUx/SMImMfTc1RF8FPMzyYj5GEcSznD+Ydj+u1Ms1r7CJNBeQoh
s6+3hkG+/bBYkmzmADxBHftP4VQccwSjohwK3wHLDHvzwjiK2GKi/QwiFl2ojfC3TtUxx2XiM2EN
UPyJ0W9ZOcwRZGX5CezmkrA3rSMlRWvf5qk5V7Jlo/i7SQI1XjgRPBkJmuhdTy3Yt3LpOByRL70m
d83zTY1tOFU2AR2pcEba8AD4jG8enjG0v95VnyJNIBmJVbOq4D4aiLSKUEpMmGw+pxSPfRb8Lmgt
xpgwTxoSy/MO4BkVg4CnYMuNRk069ZBISFCAK1OQ/VdB630XLDMekk1Q4pNC8qiviZGwVzyx9SjR
L5DLPrTdLZtq29NCUncnEkTi+gMsyAISy8Y/sBzv1pPnN2qce9QsuNl82AFOgpVyDHSwQr7wpjMM
smmMeJE0L7CTtDTO4SUyQncmeJY0dqEa/fcb+ecU4Q9XG24GHVfMlKnjKLetPKdUEP1CVWT7FN+o
FvgNMdC4BnE7kecubzudfopdIZNL1y02Wo5ZqFYl1+/JaGCjA6YdMQnFGoY+BwS7KgTb75N5b5/5
MRIehtoiBheMfcmzh+qppHlHthFgv0yiTs6trD4FS1VpCe2QDx3JEkEPwaXsqkOZvWJX3AWe2+66
5LhSR6GcjBMVkgEOAwH7E3Y7eO9XqcQ9fybFXsMM02taJwQHFgzvwaasfO4pUksaz2PiKrdFIKkZ
u+7aQ98u5OEYggW+Oxp+VgXf2LU8w/qjQnnjcEut0eGhe5zh2CBQ49e6kfnojdErVhhHcyIs7zyc
aJaOcFupkrgDPRh4EqVkZlivm7uJ6GcsTqqLzNoj8hTpLlucsd1YYIqeTE+IDh7LlLG7diRDt0v2
90SsONtTDCsq+0VRDVyjDIqnPef89eE1beFZHNRAyxhJ7aIYNu0N2c84uqVTaynL6WQZKfPmNNRz
Uwn4chnt1MKWI5t1+ty9Lk22Q4Id0X7UPjzLK1FvyqXQLHY75F3rzKtATVOY6+5EDWytPbpvq5MD
EEn3DDKG/BToYkkNjxZJo41soHRDqcYQoR9Gbg5ONXzQOcozdAwh2amlTFXTBwYiT7oDwL849fmD
3yxYyzPmmpHubVYJtnOtjkyFESg7w+VakdAcxXPHlgNXqRItG8L2nrF+4B1d39NMEeQJvGXRrqIr
FbOI/KD09Hf7hpzCQPtRZFIjlXGEYbEuKDaryc0P9elLeAvUtU18QhcSVZESJ03CEDyJjxkSYAC3
m2PW+ddd4mHy5zD15aO39uJNWLChNRDyjhudQEphdCJYthMQphCMbUsVXv2w0WCRGiQseV9PdON6
Iw3hjbv5w9onaG1G5395Bd9ZmnDewmC1CIJ1kVBGtdrM9mtVY2SNLYP8cUza/siHFCtZhIQ0oS7S
5g7xCZK+LyQlCqw9hK4k3QAbHMoDDATnk19WaECVkHFKZvFY60LRSWzQDZyqst5Pv8PV9lS3vGYR
vl1ioYVHQeqeqQCmIswXEcu3EvA3Cv/5CHUX+418VOaxlv6iELYZvT3fFBFgx2xsmjlYCDJcem+0
Yrs/935A4PJtiEut3XTYwgzR9kpQEIIcYOCqKFSrCVDPgxjEGcUIUrOKZiZeHXkBMROJNPdw5B4G
H1BVCAzoPhoNX9v7KMzsQuhoRZNdaNiIGwCDE78q84xsntBiLcrMFF9AJ2OIXdRvFHZ3bkHyGdkA
U6xjuX9bzlUdQpSEg5I6epc0sU4OoaLfIuwyvhaabTLn5ejaZPTJYDwpT0xOKsGZ6P0ej/SpmPPQ
8NPXy+fmR+kS0TjMvTQqRjEMcWnBPS2LiAddzMnKwCpZiN8tNpCgEpEoIwgOE4jejuWJJaAGXkEY
kMFaYVKY06cGLCnr1LCxb+Yb/fWJTPL2u2vWlc08kDHZIo2Bjaxc4nAQt3RVqm4k2jVaEmtd+AWv
ZmWbIo6R7rF0k50Zqz/3u8Pm9QbjutwYuHnseuQZkUjc+gm/hpMV7q0AM/rXdr1pPKR5eOqG+YNA
zf1VfqE6MKzFxwdNt3qQnCUHbXNp8yi14tAHYMImdeYZtVScfLBgb3Gi/2EEH3WW824TUTd4jI2y
cnbf+YQw/v6EOBUKTmKRbLS4RcBp5X5+jGa3Mplwtl+ta04nBQACmYEUe79BaTRLnfPK2CZ8wuiI
g7ElKpBDyYHRc8ZspARrg8HqW5TzWJxs5tbd0A5ftr9A/+4q29wqjdLJE2rJLLw7P0OCer1Ak2h3
u4shKkaJquDnzwOLCgeZUVM3AD18eougfpWY9jLJqbJAHGo/JqY0JRKI+I06UwU7zv4vW28vRYV+
gU6M/Pj55UW83VYDyPHCukxVcoK+2xxruL1SctEWcm13YEdSqlFez/0iDs5r63XYSuUtVN4W5Qmj
fqpR50XOeVLZyxHbfyKbSt6iYxRAaoWtHLg2V4rRCxiANRyhTLwbANoMsnz7RlcdpvlMMKhgiEiv
RAeey6KTCAWHJuAMSDbVilUBYbtVgsU+06a721XfCOFMGt6u+Ua3i1tP+HXVqdV/9V54yatuargI
acyR9VRJCcW5ydAkRepROQl8vQN3THGrHtgdEEdkkc8NbdThYsY8IK5ib5uSmQ06k50PXBUxmTdY
rbBwnbs91yTX9TvpxjMjeE40Kl/bLyul7zkYfHOiHF3gIg429kpxWr1Gs4QKpEh1drcBnrElKDtg
/WuOgDYQs9pJt/jsfm3H1hgxAMwi9veKxfChSnBR2Eeiat1isls30gbQ8DUmg9j21EqT0EQ4kXBU
ATyBO45u/QrQ4hyMYxf2o4OZ1rLQ6xMbUfP6fbjq6FA+46h6O+YVTMqhWKnetI+LPw+jxic4Gv19
C1RI1yluBXVoIHgKfsbvZMJQhh265wApglHFONhb6PorB8oZaZRJJ1CjK8jbml7qwi99RdsjOSRH
9jrf32XkpdUOCmC7b5xPQdTnKRTqnu9IOA883ZL+FjeA6eM01k9crJDqLsuTZopMj5BgSq1hkbHl
t45t54sOAsuLoIDFC43zBA9bueY+LD+kR/YVAQ8+NFy3+hzFQrtwPlFs3bafaL6B6LunOWGDh7D9
ZV5GgKVxfoyqEL3vR+L0nTpDx7jrGa/rWJBawSOn0XWnc9Kik+tPilzPO4rC6Ve1zi0C6iPG5zrt
vgpgv7wmpDGFFbBXTRtzTuxuVdjG9ufjgi35Oe98HHqMz3uauDNNAIxa8lUSYfX3PRRy93LWrObW
7yQnIwyxCpykd5d7HIhQtLPVxhXEmHCh7oRX0+p1jbdY3eJZii0kAacVqLba4/pZdsvdxikh98IO
7opg1waCw6BCcvmC3R3SBqsIbWStBROYjUlV7uMHojPajHR7b4II4hgNZeRyuhbFDwmKg0VG56VY
JHoa+Ml/I5+KA0mbyjB/4JrghpBkB6OgODfboqzaZrm9QvBWnGTjxZ1mb01D40kFWZNGXpCmAudw
QP778bmHPTdjDGeGSuGtS7zAhfvvtdvMy5hv8mxa3Ymlsw6LHpMovb0FvBRsEU/gIKFnbaYUGPYe
VRhcEOIe/hzYyJCtJK9xcKu43UKGbYIXARHPUy3kpKxUBDhvL2Rx0xbTrlywR2tOb9PCGFbeYt1f
cJ1rsjHvOqCJ3DL2gZpQ85u+f/muKysDUlGNwMcqF2FbIRzbqipCx0YsyUT6AeCadzTYjr5lbjnc
CI665T6AaoI56TWTo0rptidrY1kZZo90cpFfd591yDFq6KK2ABdVVZDZfRJZJiQad4CHnKm8fMO9
a4+P3VJabxFj9ovkh8ChNE4J1iDlDOEdcZ/Jwj+4nKdwLggJizuupDi2KpiSKbaITpvZDiwIeD+o
0VWsD9Jr8mDruNfAoKhV7+tqIG/qGk4xN0033MZRroUWWSu7cqXK0KKUDlRvaQRrzxQXDeE3eT9X
UHG0WZuTwHNZshiWysb7SEZ/6yAJMXQapuZo+EUw6dJA8b7tl1Py1WjovMsH9nLe1lFKJPNbYdpH
j6ZV3+DQlS7pu67vzg4faWRp/nFqzi+s+STOpmnwGBukhiNq2MNJg4RYMJ0cSMPcN2lpebXoLZBo
oF8Wl5qTUVT9n9QwGxNtuUAVlOhvwSgCP4iV+O/bAXqvi1DhS7GbpAkazOk4uo/9qHiALGbzyXe4
2q14XHJbP6auYz9QosmIjBnkyqmKv2pePQ5WK5+8JhUpSsvmxy7KhhEUunrvc3OwNbXSYwzyQ7cj
UrwB/BGqjhRGZ0jLm7TeBvagvK4Qj9R73VRdJOV8E04u4gAcklYb/CM2wkC9vE40Sru+J3tBhzQh
Ye2XcROvC/X4EjlneNZjfuH8op3T7qR4hO4hmKvjXxLRO5CQSA7dFa3D948MvCREykdXZe5ErP69
AmlM5UPjZ20A4ffJVxsgnIZCQqRfs2sXbccl68pbeS/zBcQjPm0X88crJjhV6gOAA5zKi7TjlPel
D/DQBYYpRAjKLHv1ZlV4nad+3UzamoWJoNyLgFTGJX0PaRw11YKhFifFUVtE1L245G4ZnM8lK/OR
+Bfhy3Fk8CJVnQLGB/8q+UMn0rV7r7H8hSjDLFbP/2g4dmVVfn8n4q7yH4fJFmSwZwPCymJUDYbL
+mpKp6xAkGjgPWaMljR/J+eXQkk9Xt36SRMEqtHJ49JqyxWStdl6XC/b90JGkw9jyfsqW9pBFdQt
a1gKRE0XI4+N97mnIds2oux0PyXVyASItTs563SF//4lD5uWf627f/zJuFcg+HQxvV8fFQDr3MBh
WnVtwTM5ns7QiTgoElL3IGis5Tyh1xlmMCKWQM+6tPLo0EuYcT7tE1VmaEVHTJTp/EWdMLjyoJ1F
D92+0EY9COia5H8TZxO/jG8DgTU9xjMkOPGOdWT9IIFcggkJir8WL1d9qQlKRXRXQc8VYBXEZUud
LFZY7xoKwlJqoHMheq5pymQycOxQtl1UyO/BieQO/9UserzWsAAU4PZt+AxIjFXk37JW23PZc/YY
e15oAyL+5mNnhwoTmqoXgVRiZNWn5eEpPxnfuDkbRplWwQfCrLByKwCZBoe0vmB854qGAwNYxKtt
Uk97O9bGU5R2VYzXxsGkSelFGrS1mUtufDMcSyA7j7n+8tBKIXcLxXAzhgDza/fSRu8croE3a4Z8
fhWZeUsyrQCgtCU7gPWot0M969LlrxKEBi+WEq1B+/mIcCQ6Opx9VDKa/UHfpxt6oM6kOlHhsNW8
BWIYHwsEt94BXVTprTEJrEBY7j/PrGPNsIJNqTx6Su1JB6cTST2EjfLnQHHU1ZJjF6hdMOXm51kF
LAziJEjaTByFfFC/19Brw4coXC0kUb9pGfSIMtBm0uw6fzSxiyq3cBXWuRIrrQFHiM2IMw3chFQX
gs9Qa4mIp6aLpIhVBIzDG6jVWxHoZjRUitoDNFXVSXW7ktG6OAuOr6vItXqJPhxygOGLRtE6T8W8
JGq8x5V8BJ+V/Rhiz1PPi1z/4P8i9YCwEdaN0++/MJbjPXWe7NU/QHGZD2C4/MdHncXydoHc8FQg
QXBL2bot3TCT6jB33td7afvB8z/6vNnVFFqb1KdTFYaC/7jpKsqtvSCGQUfjEOLnswsb6Wuy8NwJ
HHYNmexKyJ7uw8EdudceBu4hxVsx7cnVjivA0lNz3++Z3rjxnW+7kMGQOUhdJB2IhftpBv26FtpN
GS7F6I+66YlV/xKbBAXsvpZxE85UVuL82Awjx4TEpPSfm9WveD3fHpmWz60NABxzEHKU8fPiqUT+
MP8ju+ta0r3GdDG4zVWBozP7lo7gHe0vhXloXvcit4w7OlbP0ktcTat18Gi+I17/FDia0WxU7ktN
C9PlgDxuzFVP07BTmwybBBttTyy+5iwcCv5R2Z1znko7Y4JodiYCxxIYkrPDX2ivjlvACd32dEJe
OBSlaZgnqB4w/SqrTySiIUyzF/kxoh/3Mu5nHtoDyp/IhkACuEq48G4m5hlIhANjcv11CM5X5jZu
DjCQ7oG9TObRBjiy+wX7TYlGT/CylWlXQiBCwcF7EarRpnDsPYARZw8ObRcVZ4U1jRyvPJItU9NQ
YoawQugk6PzooyC2bLzshRHIGEESEsaPTLtAQZpxlyI8AW/L7M9ir0yZMka88j0K7zejQn3qyKm5
FJdX6S5HK5Uuy7j61idzolPXNvpC6UF7riTSAvhclBvHlEvVNvu6a+vRrP0qPDCr6aVv2AIyw8vV
tmYNE9Cs0vYR9Je3Dj2+tZRhXGRVo4zFu8llebzOWObPdL7yNmrXNp1HLC8FdYPDpT2z7he6kpz+
b9l24v56Dvke7YAK7pIyLfaySxAdKezk1z5lExxxsHClg3yte3IPjYF4P0x3YPHCyGbnQwtkpHQ0
czdnQcmV9GaJMs1dv52DPq6gyeauoZDSN/VhpSQ/jiZEFASjhHwS+gdvlRPqDNlzRacgpcu8hrkT
VeX11Ev2+DhiVAjWXtjjtMC+h9MT/wS7PkrhOAiMRuM+r9dp5XNgtrrpNJWnI/OSttvPo8HLBzW7
JjgNyON4Gwf0fIdMs4W32QXHug8eK2MMdIp3d+gAMbJO15euW9O9mqbRqhYp/UAv+8sMzppHs0Oe
QKAYkKjEbxWdsC92+kF/4e+4zKhji3c59zRDH0R5srtWxFnwQHRfpj6TkwYQ8MHDlr/+p17TtIzI
8KncCl54jEtIOUnII/uUlPkGn/BJRjSGdOa7ZdvcF4NeQfWy5+ysIKwj8Ji/mDGGrSLwxq2TIycr
UPeUIC3NVsTs7pBhMonK+vJglZfUX35LUB8mqz4gTeUPAEZc+zZl8xsNozGsUGE45Y7i1wQJOnBC
0+NzvgdQbh22geDPRz30f+TUtsM6zig51uTShYFiSZMOWrueqNlwiHkD+TbVkR8IJmHR5/eXorSm
ihntRqJtF5s+PyF+M7X0NSTQRI1e1ZN35I20FkuA13BJMfBvKU8k/IDpcs6uWaPfr8ZKstIRjNLS
fvCkw+6OU9FhdGDxAqRfCYrajo9CH8QbD4KjiwBga/8FCO/ZDJoVwmgKWNt4JgHWalC5+c8ClXiX
YaKiBnsF2bKU/E4ZqdOLuFYRKStrGV8UuplHj2z/TqO06jeo/SvaM3SD9yz04m0GMQpztpXu1Gp4
i7WB/SGlj7QwZ4GiXodaQmilsUiX8zvFlnto31vA6VMm2v3Ld6JFPJT+nCXJb4ftBDb+7dZLJzIa
kVeEFlLG0gtxlykHzZwYn0eIhLabBHsQcRUQGp7BjnEb3NKWWr2gJ7Tl0DhanYEPgcf2V5hxmpUX
TNpvwc9ubAy5WCn5nl1G9UXKUAHV+IAHTbZEapRn58rgFhofuojt8oBBSKwkYrmXJmi3NtSgnoH3
uj1aZhmUtWqoDmnzrrgj9rbfrSTQmFIO8sn4YZak+SAvB2lbptx+fGRLNOjHc2e7tNwFCCEz4FTt
yfkntLNOb5gWHp0p1PqEkZzT3U1nt8GHErSa5F0erqCNcSvlv2CYcesKPSplaiShI4d87To7XC6Z
Y/iPsdvjyJe6Vdz7gB7+XuerBkOMf+jEqq6DbgTP+3LZpWs3LnrHVcMXzKPy1jE+iYWo25r+/oT8
31FGgfkzDe6fIaGpekQZW3hSPiIFVUSjRp1bNcYA69dLXErRmpDmsD1q/EaivSt7Ibo5qWjoZbPp
bCE6f8xQis+kcPP2tW0Nv9LVTEGD0QWvP7gYyb8n30VmO/lqKrn3mlK+MCK1bUXzNRPAnmSU54NM
LbdOYGnkmpPdImRLSjJqBD2Vkzqb+xSDV2IJgOALH/oYwnoc3En+22B5Qkfofaq/qjwf5euqaOfs
dip4gZ1vA0QCNYshc5B4c9arCA+Tb8lM0m6bm0dDkkdaaLZWZpNzUZ/M9LYKhzC450gfmwq+1c0/
FV/FJl9PdsRvIbrMFZr9Fyq+s3rOxPcJqHxNgjYQT9YsXsP7oUR+ALJSg7GsfYra5qEkm1vapyhM
TRu6dHw+sO0DFMzagQ87L08SKECyBaUhsQePqIFi1HKcCrzTwwmFjPY1RV/HwAFHLwtl26i9+BJM
ULtNsBLS1DumMLnu2kcWSZCPpFgE/H0WF2D3VO+rhBPcCqn+1Bo2U4jLrxpGSpZorpUrdiYNQEQX
AWLDTMDFrzVfoxxS2HXMARb8qofJp4u0w1ZZMJR9RFsC2dtX77P2nyhUXe/TR9j2BQLkjIfe1WVB
7erOUW3DlrDfz2M6NxDzC23sKieT7jGoD6iTGclntsSvXKvBa0Payzh4PVyspjzBXXh6IQlfmEvr
aTLpq5X0qsrVtWtTiC92+OsLPgLXNHmCHpBbtfPRQB1O9ARbXbEZQtBmKVjQoNYc186e9MYKzIGm
JRfv9q0d1F6ih3IW7CjJV50F1xokMeFyacJrMm3VCWqwE1aUwQliSROs7Nn4R5+vBzmNMBpR38uM
gRpnu6EG+UkYQKny6eeMHKtJoCBaCaSCLhfN70oHDKtWzhiu1G3UlsvAXtr4XLT5r/VFqBr9t0wv
Jhd6Q/p5qRt5Dt5Zxd3KQKXcFzVBYJ0eqgUc/OKlgcxcUuVYEIDTM9APcMvFB7MNIdX1J6XqZQz1
14aH9vQBFQH70r2ea2k4GFh72yUJB9DrX9dYWXF5jIWxYl34Sf3coFPOByfh7iMSAyYCW1oBlimD
nJ+amxEZXajAk11C1aJRGNcPcOiMEu0ZNMIbAeSDEgTTSdWIrjQth4xBT0DvJLdObBJ5LjULgqv5
okd4lbf79roygH39NqLBAw0i32SDKgAubrSpy34lFgepBE5I+PLpE//wKgEoUG/J0vm0Ujrl/sbM
BO0cddNnPVqq5JKKuoUxkis/RUqNf5VnygL0wu2pecal3WxgrsJomJLa+RjkMWSzYYGcdwO2Odi4
QQw0kCbIT1zZzNWFWuSMmak+fUhwdqP6IJqAbwkYO9OdAv9HzrJjM7sVh4bWZiRSlS/kXFzLKlhw
ztQaJx6IQTkK4jtKFQI4w085fVKVs9vMTex4NqbLwRJCbZ3nkEiiI9EQju+BiY8f7aSkaz5RX8F+
NZ7bVT0JA5UEeurClXGPpbBsIjE9+x1yknL2xxrrwjfiQBeO74B4RJ4GJf6JS/7lxviBZsi2P/NN
rlmL4S+0c00Pmv9kFKlp04Igup5OxmZ7kJZOkBFTu3KOG2w5vJDK3Qt/mnCBuhsNNUGlCSdzUUGo
LZxIOomdzac66e8vR5evTyCTFm6sAuYdYykscGdmxitDKGkYdleq1adowbbugF7s3SzFn7g/flsj
OPKBFR4J3HuR/8Qb8Lx4uHIxgZHMau30ayqszitmpeX+eA5lNSaBw0gQ6dm0APWlysLojJnBZuNZ
qryenIEK4BQeO3vyEzMw9DJGPNqxPKmQV1DeAYN+W2cOFnMFH10+oBo1v7bSIG8kUV5dBzFKfcPn
5YcTeCwwswkL6bE+glk1AhXrNv1UI3tO3qX/LSaSJOFlh811AU6zP5MB7ygU+iNNSqT9arrPXh/m
xId4njEQqHgcYKpL79jVr5NajfdmLJjs8JhMowDJZ8ABJ8/cO7ad5yV2FYtKtRJsDkujnaPbBGkQ
TkAQYfuos06I1XTmyx7rHBIFLpU5IS3/SVYtt/RxCskUkvwVdNuNWxojbbDDn94mQItj2+Rjdz85
J4Slb2XnTaszTJPEQm7LeObqKdAfT5ovIyzJs9EpL9o1/bnffv3X5tOfck+D+7Kjs5gSV4zK+ixk
11i1vqe7aQa+Y/OmeZKgNvgdb9bMKparHOaDFaMAMGevrNrAl3fL5uAsqVeUSbF5fneEf8qJd0j1
GXw5KEzsevs8BnTl0FLi/UtqjWX/Nnrwh9XyadDtZH/CT0/n/nKx00uktaned1pLSsoyLHTWj1NQ
SFFfPnH3zFjjn0IJFb0xtN38kWQgjpYlqqHKX8yAlMq8sthj1j3vTkfKByU1m4BjCGC2ULZ/+0fq
tZl0fAfknh6w8bkJHyNJn//hyOyKmF9NBxDtjyH36wEJbp9pbA+zNQ8q367kjn0izYrivLz0OVGm
FEi0C+f25FcK6kfMTjWbSQSJMggKyK1Qd8FDBLQirgBNc50ub/CJOHABBCSC1qylZXuXE8kEQYdy
A2Pk2nMhH1v1YQtuQo7BPn/T7eiNf3aFVQF1/6k3BO1eJbvbOqOUrVqLikU+vKf/GWNyBADchrcL
PFg3bWoK5fSiHhDqY8r00TzyAd7brBvnaYSqGBDqk1sUx2KZuzNax7GFceWOy0ZKEhG5X3Sp1tET
rLKK6abPH2z8YafvuzRlYy+mo9cw2jmGygYvUfpVAjdA6j3WIcc505mFfynun8FZ+JugKk0KFGvM
D4SiHWYyOuXdZaFbZbl0xokIJVPSmY59XAYIgP9pcD2Z50b8AEyBf1+0LlZSURhwXe0eW4ACsQL6
wpChV7tEidPCS3IeRz1mBAnuBFGnSNLRpX6Qr72hfCJnriGrM2XIgi7Ntas+fsO+sdjiJCCfC7FZ
iZjmFnK1PutdVlmpN57kl3m2B44k7kbi0tqNYRG/sMiu1xGsTn3VuuDEkl5V0/Qn8LatsIgUqxQ9
1TsTtid2T+QFnAcfdQxFuUynvmKpuFA9cFc9y+TWYDdqJBwLJ0SMxGGd5yrTn/u6lOWFDaHqc1w+
IL5QrRzXZtLPrbmDoG6+kRJqIsJ3f2r14RPnqcwr6/27jI5ZFjorwYMBeNRJ3gDkDSPVRm17yk43
djCuphXPwX8qFD8dYMwP1EO9oOnKui8og79jWBaETFwWcoMz1gStWwfZP71Hkp4BqZDR+KPJl4nx
jm3Y4OoPQGZG/iSv+wMpWRsAAdEqQL1devimwcuMHiK06HVpkpq4xBUbtkBOTtKinSNOTEWdRcv/
n/9QfBgZMRsqcDeVhRIXCZ+XVVtpXccUPAliSG2HgPTtukGE3J0ifXLZFKcqHKxyK9MNUWmO3AZw
GIVYFm4kgyTODksiLavejU6eaTk53DHU4im8uGi+BB3QpdQpMVwqiM78IO3tOuM/+51hdSd+xS0M
1M/LTFSAL2JJa1txhH4txUB1NjWs9x5i2C+tAJLAIjYKJTFvsgEYFPUa8yDuqQoJ7s9GPP/h04Ut
epBfMlJ3621UE7MXIuXw/ud82h5yg52iGKnKt+25AcM7w8Qfk5CTLgCMgP3bC1y2HV/qtpVbzoth
bejjdgNV5EMusp/uzS6frGjYZazGT6V47Nwn70cc78CJ385KywB82kNiB/vxWkuiFQlGVri/wnyp
nq9Bj3BPGBiR2U4vDPqkEFtL/4n192V+OA7k8MY7GZLKr6Z/fU/Cy/hx4Bt+Kaulha+vgIxZnexX
XIG4tJisIq0r1zHOyPozqqAYhaF+lF91Cja4RNXUY6iahXDAwD9Nj57OoL97r2m5RBHlS4rgrkqJ
hTzw77762Wm3vL/RJg5w7bmfRV8rgIPtEOEADwSwO6puOWRWDyU4lA7WKrCzu1FE3/S3Z353stQV
ynyfVjbJmSm60Ls0qDxVvHQy3VV9D/NaQgNuxaCtpKJRqckFrtu6vc8nL5EvvVgTRN5mqHSeEoy8
oQ8hQizMAydOmdXsZku0y/Zg/o8IOocINscbNI3Ksh1+tlpY7mHIbOzUfRC/OwDt+9JtY9QGAAVv
K47cy4kPjSx2WiR4eymdXXfmPUBOILEs1GJnTBE+ezBUpgWR+vrbPLErYTx6NXdy7uDc1VcAg66E
kp3u3RAB0iXTSKav1gHO65JxpwMdZ8sIzSQezb/lL8O89cs55iZYsz/0Zua3j0ATfigX7NazQTiN
9Y4IAJhEDeaTFD6yOiLw3abZujNrgRcRfXzoctbyDlFwlO0Bhmb29YCRG+YqI5uPvoz4AtDGM+zg
MVe/NTifY7ZHrVu4tvOQWvOm7exALDBTQgiMfYbu09QEj0I86MscBM745rDFqHqrr6GFDKXzqkAr
D64d1x2KNAVblBSvLJglui62KtM3O7g1BDqE5YQRuWedQ6K7YY6uVg3aneOfg13C5xeFYQSrMfe9
Fj35XDSRBCzI55nD0D9f6fzuxf5A3o482lfSS4NNiXimBAlu6j2A/D9TKU15jCwkcl4p8zv5tpzp
gva7qjWolWuZPGSfqANqb0+DKK4hZYyyU5xdXXYrie1AIFpVm4dMhVWjED+tH6uEERQcjbZ8HUdg
BLFy/yzhaeyzrkCFNzgswLBVFfv0I0pAtIKpmDIUCvi6isR1Q3q7CgkWOzKI1NEPQZXdpxgke0sF
auqGaOzP0bFl0+MAOEvbEocHsSmzgXZfga+xLA+0rJl/v+yAxI7IJIyGqGJo/e25Gmc5kITxAV4O
k7rbJHjLutJP/MN9PLSu3jTjI/5iZSoCtuJUWnIrOhsLyG/d6snLvFz6lxT46Gef9h4RfksuT9JU
aubcyy2lw7a1PjRRGeTfpqtAlFphLstHYpcMcJA6WqcC5AMkzjVRZRK6Ei/R2TB3uJmokShgG7sm
hgu91iwNZUqmMqgNm503Xpp1uh9cPQIxMggXRus2ySOIjWe5P61N2N9JlL1lIeWrg18lSLVDDxcY
yKGwx2PllLnsvKiX9HZ/8UH5tPfNTBuD0H/j4hDLKhI6SBfftK+Oj8V9fGCZwiwNq89FAtteM529
P/cLwCyJeTxeaO31X06lCB2nWSYoUT0rIzZqATg6Qfv3UIRUiXhoCoMNh6PfYsy+v24GXQuitP9f
LErVtp1wC382cUCgePwY7sTb5HklpVaj/v0uR9W+j/ZtKNwXVckRmrBPEFK+SbyFhrbSn97yffw/
xbad4CFAyKYMsdUT3EMZhybtaOIkKhEA9Ll+zHwUwMVAz8Tf6SrTtkynYIO50myCXAfGmbXuWPBU
SxTJ1Qi91zyGrr1h446KKeAzWv3lmknZ7DFFZwL4xZNyU1c3GKW/jGqErP9IAJUUkKjv37mPzz1E
HkSZSEB/9PQcmJyNGnm/WZ4m2Ld0k0wHCobBHjzGa5ivSg6h4zqArbHK72OGzMglOCM9ehmrjjGe
dkEQWkZ5fUqC9Sf3xPYfntT+gFKvAJxgQUESLKhZSd7hmpMJ+2TuvW31P69oe6knIy2ntGizwnpb
ogiaFh+bBj5zIe/O69g44ReMPvbvsGK1f81R2Vh0hqKDGVMtEDI/SPg/tMxCBOr9VCtp+9aCpulx
KbaZgT9Aa5ewIzIcYRqvs/kJJdUL5cZSy7FpW3fJxNe3nSfgTs+dwAgA8vO1eh+MvzthVIEEkxnb
Woof04Wtibsmf+c1HAyenv4owSLj0q/A0Gn6K/TvorRzON0LTyyR5TTHnWmXpiXVAYS8HDuKjops
9akMjrbNFkIp/Or/QffpkY4xZhdm8CuVpznttiXHi6seBkQk/qGH0sJhTsctXQ3yKNQjvsevTPBE
Zp0qQmA34b8HGPYrj8ui+dNrKO3rZQwpe7xq0wFXMmQoy6koZc+syK8mSzKNb9H/VumwN8Hiy+sT
2UmWDXmvh9GvfYA7KMAV0IDR3ULwKzlH+mQJeyiN+F1rNEOafidi8DIB7xvSptVnf8Dmkn9lAsmE
nTUWyVS1WlUaCgtzP9dMzKixdux8W0kNwxmdFJ4amG0dnghING0NEl/D6W8Ng5NEbY0NsfS5B6aH
ROwrHLTRatAmfHSh/SndYfK/atbgHLu+zw+xOeD9Qo/m9IQIVg+r9qbp5XYEx1gJnkSSpRIy69Bi
LAMnQDfUC3XhuPaE8d2BDiOk2BnkLkHWcQ6fwCkMEA052ImmZEu0vvCVDBT8yFVhxC4ZNMZlC42A
19ju2mdOglYmIJVbncmcuCQAAXhcX2y5hJeSwoqNuGOK5OjuklkkWqhb2QCNuYyKSEkkcpFPZ8XM
QIri5Qp3lJd+ZyIIOqA4wonEan2niOgkKDE2HFynbS5sAAYWlufpmJW7xdIrlXca9J0hDoVBfrpy
3GUQld0b+WFGIBl8aRCojNllyycGDh+S4FLLF+UPv3BY3rRNKclusAz0RQz0UgaEpBs1nph3THp9
b8BZClnA7mIP65FnEmnSHJpylGN9AH6KCToenye38TzSA5UcJLJUlY6A8CYXJn6V8znmZsnhnz01
/aec4axQr9eS0A4Vyg42MP8bi4eMCM/4qVIQwFHRN4M+cENc4LrA6PE9NRKOVQVkCjZrj6RQn5HL
h9nPSl7Ixe5ndOQPejVSAJL2Hd9fae93r0dsW3Yg3zsb65TSgM7lKrxNSCJxWBT86gluTpCdKQGo
QPI8hkrncRO/dUneIuPBKpRDLLGq75IO4GUwSHbJsTOFtQK9Mwu1VaAgFz7AQ+mCt0ktOcrN4ctG
pS789S/xh84Y/I+cmjDUZh5LzEwvC9ZBtYpropaAgWGlbAxiDS/qWLL+qWBJGMqBJNQtk4gCBpsa
5LvQYHY+6qroKLlhBm7rSbFj4ZQzthjWewLh6xxSLa4KEGokvd5ZNSq2lsqGcf1d9dNmGf9vV5kY
sttJEjlaZrJ4DZHO44hZOZEcBk7z8U7JNX2fEWor1IRa3IgeymHzftpxhCbyu2Xhc++mNzih0S4Q
C5uvBYRA1tuurAVroRaHELxG1vqqptnQ/J894H1p/aMSJDrYaQM2xo3TrqNOKRrVTqhV8/VqMo/T
iWdmW0ZZRgWEvzc5X2KafRnKrLlNFUiklupCZv50Um+JLfh49TfTjQ0ee3e/8xrP5VIeHp+qLlTk
PXxuJV1hc04RFcUyrNK+1Nhp798Gtoj/afrBneLJLggw+i2/oC1qiGAdQBTaIVHEZ+dPTCmYiuBo
tL3vUieVFYXELAmdlsosLWlYrpIVXP+49Ld6x0NnoaPQvOe7XYniuXiCmnlnDLd20Wo6quuX4bRp
rf5Du5zsbt06xba26vaia1x0TY2KOTddpFs9fQb1mvYDtbrq8r1vyOfisuXr3R5ydiiZEODSdgdT
NZKhtfs/BuI58pzDziVhoWaZu6Lj4C2cWLXpIapdUgLIagl9PiyHqjVQAtYKG8wJH/q9tkbm5aAX
s2VHFzEtQ+34uhODLxPfv45pd5mvBnkyPzVDB4wRCVve0sTA11jMIR+EwjazAiuKzLMvAIApRUly
az+wxi+sxfrRuFcw90HMgqsUV9atPCUMeR+FMCioZKRYKCB0y1rIQAien7cuSy/CbnRN6vU6TPbT
+1/pEBGrAvuiocZeQql7s3RAsNQTAbbY4hEJdC3fdksJSGBLpvWhsrohzJKszEZNlqr5ciWYQfcJ
ODXVe0E+W1sxHvCvBhR+/aG35zeVArRuo3z2i2Kt6O0KLcj09UCfilv3iubeixA4WfEuR+XTuYvm
mJw6ZaVMaS9Pnv8T9UP25kXmASjLesi+NxKhWrYZfpgEMUMa7EzIKD6yHlNAGaVbHielsXyuJ3mn
MWHFxafd3gsyc2IVF840MskcLWYEoBnpCzIdOpUL6RK3Uv411zQjU6AuEz91ev6ZUF25+mQan3zG
ueZ05EoKYVz7FrIqduB/RBu+p/NYtazUG8b5S6FbYVRAZXmA2I1O/nI7t9pcntsL8JoIVuf+15vl
prmG5pgULoZixUO4Ao3Ro+m2n0DaDOBSX/9UNCBves4B644nwa/uzrAegoszwhrqcpNsEVfT+vgc
RkIoJghtUP4Hwm2+yKVegKxcHDY6uAC6jsUSUtexPA2jeauIBQyupHy9oPHwl2hnk73op8AWiROP
58t5a08kj3CfP+oUZhZ73Da4gPX4rb86cCB66dQ9jJX1UNoIDk5NUtiBVS07s1q9ufvvBAt9tvUL
1KY0Edbm8/NYIZeZ/mcEHad/Noi/KS9pYe0jIfqDuDwRu3Mnv8jFvEB5rZ7SFOdVeqgtSEsAArYF
WKlqOkjw4tKW9aHGaA/gjii0cHYi0RBC8k3Yb9DGXoE8PwH7naUarxdTJZuWvendT2G2VP+k2Nyk
1WVNLBM/Rexzxh86FpIJbT+s/sILZhlgBE9nl2IwmJd2XaJ8SRXJ9x/8wHFwLCx9MnvFhtLIh7Mm
PGu7OU0iUh4hmwu6U6Z6VLRv1I8UZEyPCdhsM1Jfs8EnsjstozvOR6E0iK+RzNoVWNiPyD2rEkzq
BhEiDmxsV/BKOebPPXUtFQs58zaWjKQUKNVlNyRUr6XEk7SHlcDAx22NnybWXJzycGpcf+kyreSw
nBd8VvO3dF9b0eyM7cA9oKI57YZCmieV4mwN7ky/6YsuNa9OvEliwfKSm8mhoFgjWCcRPwFJqSSi
aHV2fUzuAdLTbZZNzKO09lCZz/uCXuwxOqjmknrdrw1Yc+WuP8PjvkhLmQpCirrUHnP//+cNyfCx
+cpI8syoE1QygLcE88rGWhmd8CXyjOeoSILMhebXfKol862+mbs+tvuKL1cyWGOaapfY94ThQPkG
hu8i1ZLMUkusJ/aSKqEsyLXTlHZuDH6jzE+Y8+c3ERkRix+KhcC5FyFM9HA0HjIovgIn/QVVLdHz
omwVCRUspUXC165EdfQ9vxy68jS5m91Xuh14UZIkWsKOY2PP0ZsX8boKSWtWx/4N00KjP8p8yRZ+
f0qIQFfvtFbUc0tzgQvJqXZtRS9A+29zNrmFsDLJDAPZJEbcy9gpuho9Uh9zXaNPlQkjDe9b9MWS
taIbIR9ux/UyQ3joY3PAs5onMweDvt2AIVIxnqnIJHZV4gCNiyB3Y/DzwSz3D1alN13HCu+DKtaN
Pk1IHUqtf+t+XQ1/8IgCgPEHjJXgGn8rfXySxq7n1fnjRh1JXW9mbGue98b7TL31yIQqVt4BGpeg
5x2BvsEAp7iWBm6vMwHGhW4QKvCNMBA5cADJkNFB9df2hOoGiNdxalvuo53a7OEXwFC3EKqNShY2
gCn7DSWNtXmbAEz0FL/jdHXsEkFeDiJhfKeF75iUzbXGC0XsrvHCf5L7K0AmbRIRt+t6nsqeSpqx
fYmj12ZVBrM8InxoDbUPqkCXVHbNW9JoeZrluAA1Z2CFDAdLDpuNv03+50Y9SPWxFy2Jvq47Is5Y
9w4X1i8lZlNANNoUW/qDKzq4hvsIuHOp6sbMfecNNIPxOVI3bD490ksFihGePDdWTGZNB3OizyQz
YhJIA+23hxTU8qPt6N/NlmZr7PHqZ99mjZmw0qNLoZNoaxiUbfgcmKM/bERy4TAuG/9EYDXo06+q
JdrZ5AJik5gQrQ+aAhsC502RocDQoc6ELc5mh/y3IrphIjISq2YCb/X0btEIfdMDX8A7CO5JMYLX
V5/VBKrIgko/WRfLwE0k/D/hiIAEwOgNO4qVcliZXEUlVG6MUiEjMxg8f8zW1f9XQCK1d7ickAOa
j0lT/hQU2pOGYFxV51/6bobgJFsygf0K5MGHNxzl78HHjaShHigjm2/U3mtQsklne1hUifkYFn9a
w51kpcNRTVlsPgUfL8UI7BoWFljzoccnKKx8AZ67aBA8GiP+YG7i/GEQSLdjNVyRjdrk9F0H2rzk
7KXz/st0bhqRXlxX4samEE09VeCmDSExsVONBhDvPc1xRfXcMCwTlzxSM1EO/T0VgrB0BJgaUUvB
VH6IbChcq96QgY4Wm1AhCw7oDNDxtPydI0Tj+B+TEazx+wQ3vYlC7H/SkBslmRXuGBqkZqCQRLts
0ccsKZEzqit1erAYkpvpemlzaNpeb/s2H3p3wR20/UmoFPnmEvAnQwQyjXmq+En7lmUwmJyGfRoy
QeyqQbtlkqK8Hrk3MVBIvAJeF95OF8nXP448xJBubkbC+wKziVqahVJawjtnfrN56VHWxg/1CIpS
VXWxCv5a7/BsxUI39XvgV+2R1NqSmgLj9sA4QAGImuy8eMdElFlGgigwFTRrfMYp7Fzd2c+yB5Ti
e2y+Ns9ahM3/i2z9O0az4th9ElO5Tr/Zfr5m0xUaISlU67PRFj4TpUmKN62/4k4uKbUDsdmFmJbg
xmKKJS+nqxZvxk5IIt2giHfFi3FGg94M2DUUvsiI7IPO7ashKUuqlQ+d0klHjuVPOf6hhxXEAqG2
DPXZu9Up/RZHxJDJq7ywnyPsPVt+H+zW3PGSkn14l4ahZ4Sfg1FJ4xzchUwtR8q/Tac3DSYHlBUc
D09Gypf71rxG9GtHPY7H0wMV0k7ctqJ+86m4SG0jiTAZd+r19Ymkw6KlGyTW87fSrJfAIDG6Ay1v
TYOsxWlxLUmSRLb7fayTSZiLJpIDIxTTj33da/Y3BNbugEDbecgbd5p5iC2e1n5Ktqe559dsgktw
Ycdo0IkZcPW/CTpFt4hFHpxFlHhFlvVyQ1G8NA/UXj4YJfWQlzGrfKub2jjG1YOhfN1Hf6h5E+RM
mr5p+t/d6fV85R5jp7EXkO1avnwIB9yTb0D1c+MVHtcc9m2hVLAVZefch/iWE07PT3EUCypExfLB
FS5ziZWpB37kpydbcI6dQQ4pqLc0/Qe/zu0UykQYY9Dw3J73XK8BrvEvlVGp0bqAgjtrrlGz8xMg
3TFtdh/WRwIWzj6giHS+bKPssl0DJai+uIMqr9/uHo8v2YAorY4ni7uKBbfvNiWLT1INRLpPGZ2V
mKiyymopj52XjWo7seXm7Tn3BV4zrQKE96ec5aE0ZGwKX0HqgvgtNJnCN7vp6Bf4GliV1JHgmVbz
1BOJTu4n7qMQjAVyj702zkPc90AoUv2O0I4fZjHDiqN0zCd4KXwemer4A/wppWmQ5g0YdHBkFt6P
5R8bU4b/Tupq3z2EgSuScps4IPRGBnvbSt5DmaqWFKYoEm/OQxOghETD56eM7l0E2Yz1yyNFn8ua
x93Fu8qRjf/WjZnqKEdRPjrrSyPT9CJZ/Qif/2GbsLDaJ5EiFnSzlyI/xYecp4lILQ3r1JrJwm3R
p+U7pOlCmHx+qkENPgzd0nlonoP5cFzvtqmB8FKh3b+xBVUQ8J3V5I/vOHO6lG+QpWSDcgC4BxQE
ocRWu38gaAObliL/OWoB5qcQ3ZLpWiRpU7lL5Azx3+ecMA7l4W+yhr+bpS60rB0+LpJsad9YixT4
ZVhhG+Ohj/pZm11WFa2PKNGEaJsj91anvvAZFaHiebvZHLxYESpGmF4qrjeX1uUTmrAjdxX3sYCX
fjHLgbLoLz3gCS8PQHNbui0xvF9fXylXHG6GW6kGx7xApXoR8mRYBw9XP0zKDPOjxkjdc3jKfD/X
YlVEUoBPSiyu1u+ZJyqLjGCBE3KG3zjKdCSKSQI9a5QocHG0+fE3ZerIDuu8cr/rgDdmQ4NHV/OV
CFL0Ar1nGGnbrfH87+4X0piXa25zEOusq3piTpTxwJCqypr/LyqRr5GJXqYsLzPTIe7jRZ0NKNgA
5Xn6ZtDBrNcFlKbcMUadneFJKHymkI6VpKdRrb+lFx1Iz5NjCUjkwX7hlIvlBrTMJLRY96aMkDgC
Xy9f2sOOOmFSC2Zjhe5Fw6JDdNvwmCPNDh3EQ6HL3uCmXOve17XXRmBvMVkP19fDHKavFIkGFEkM
dqaC0iB7XVQMs7B1MDuaduRS8aLrYu6W0buwzsuO6ixj5nRbPMPdRAPnAenBrPTBMLTeCT8Q9gFg
zq6Nt85dNhX+TmaqGDoRN1lTvPiMSByaEv3XvIt+m8I/pr/hqb+MPDtpaMo4OaKsgSNhghc9OlG1
H6KZUiYBkwLpcX0owzjR+dIG9sc8d7WUmdGC0FZRrX2aFLglJltNEQDr8RdW0YIy6DZuqowC7dzH
V7ZWtGGsSm+RwOIwDwaTlDEjpJ1UUmkpbnHfrKr0ya+09AWQNYmTqLyw5NK2FBKUBRIWwNbo84VT
KQ3jq4lGX2f6KvzTpsi3fTVhmrEUFZJorunoGyaJ8p5bt6fPtSi37QDkZTuoYqTAV7q2ZWlqre1f
B1a6O/Dzp1YWKogQqeviuc/6DPz/hsEuHjz3Uh9YJYUVTl36Flg4EHnZ2XPYUziNRYB4yNarYFFx
/6kvX9f1AGxCahIvNomuiZ2rnWvBH+j5oa/OV5qc8c+AWuQ8pyhuWrmQJEG7dX/LX6oVrlN2RvOt
o16T1UNZDCCY4pa0CgVsXB14MkPxe70UUwCF0xSLEfUyJMpa/2vz224q0VmYmU6QgMnAHWRWMsoP
oXsn5kNhfZh1fk/QSOH1OsKRNB2ELC0tdrSIvi00nhXSOwo5pFRZGQvcITLQdmz+vsOXsePwb5nc
0q2XiTcGQka7ogjvHU35CFU08tcpNiKE4S+0uwxa1SsoyGVT4U2AbcT67V95vDtw+mFPCMbOj8KV
DPUu0NSbkSxLkjFFfaebvpIAYOmxBpfAmyOHSb8HoACzme746K64i8jX27vQuqN4yo6ommXYgPfu
G92CWzPeTy689itWuAGDXNsFDPA53tHBZ+DofRci4o4xhqcz4wO8JdHTVtaPDXeEBCicfXORP/VJ
WGldQ87QJ3MmnEFzUtM6JpcvJpoeWm3uY+J9V/zFvfoeEz1N4HnmCOhM5/TPs8cDHsFL1rANGcM/
+JHxvRr2JVKWTZjMCpuuMdDWTSKKSI2EgO1c/Eb3PC14wW7W26AV2FC6cabG1Xjv/epahXeJSLhC
huG/M3QvMrDJK0YSIbzsnIx6/4CiPhDESSTJgpoYxu/dgn2N1jOK5G+SRismIk5OC8psrSuk1sHm
Ypb5mwQLebiBOacoVobbIkF9OI/hMJWbXoHldnVGDQrAd//NYR0/4WuBGOQEOoqCF682kP7Nbvm6
rUMMwhhH0qeD2dTiNvDJAtGyZcWGohhYnXEyyZQWiS6rsDCUbV4eU7RZL01unYij5cm05fS+L8oT
W8qGBItJD3DQryXtNBfITpjpDr1qAATpbbpRWERL8SntnAxMBYM67FnH25UCZ2jEoM+LH8cFnFHL
LVbji0g9hgU/Yy1O5LGkuExKfoi7ZEEkzMf+3VSqu22WRQJric8M0Dj8skV3J0Sw+Tym50DCJdtY
WSUdX0xgoXU2yi67YPBFqvCU7lFofQoUCdzrbhUxU6FPwVvNwEr+TOSZSougB0R4UcE19ek2BAgi
9nx9J7P0G2OfGUkWVhq5FdNYLaCxFBmar5T5np3JPYEavZCWPofd6t/QxijZ6xJStOyYN8Cbdp1c
Ahs5GcS3Kl7XAD0GFcmgnV/+/N8adfqUQXEuURkkDFCn2zFqytb6xkHiEo+uCsDeQzpXfrKPDUZc
Z2zCVPI0yXePGA6Nyba9092VigFldHtgE3T1BJZUk0xMfT+SUlCb355fHha8tft13jD5jJcXDvoD
MTUr3gqh+FZKTe9MfbVRHJTp3JkTaxRZrWRJCZTgBfWp04gDBYD6cRHX4Q6pQA3iGa732CmMnZp6
kWO875R3GJ5BstevOFIS8nWSbSb2IjcgUfC7UEq1TULtF6dre908URprM2pdyUFqAsf9xyI98Oif
aINAmpuwX7cMBOt86VSVn37Tc071n66Dz61IxGfs1FS3a6Gw6trMBeDwcO8VCj3f5h4pRyrM9JC2
/0U7krFfI1zPsb1EEIyJEhx7lDbcJfe+hjGwzUn/X7jvclhMOjj5aah3zDKgSwvI0VPirKoUg5MN
uKSXHkAi4O//hzInT+j3TNfZ6RwO0KaXg1hzcrYOFYIS4az+jLTZ385/+yKx3ueIJMCkgKl3w5Sx
/yi2y5ocvnKputqj8iqwurTqMSzcE3ZtrcbWhY32+KjmRKmBIHPcyqOYcdrlrCLTr2fIIRpojjhr
hr81xTcfughereUAKSPZZQsFqNrps76EM5aTpwqkf3jlzlTE2U6YZN/muyNm+bAIeho73hC+dlyS
a89IwXqQaE6WdEPOVKBRT+6Rw2r2VuiN7AmBFtg0TPeqNn4wHJ3uxosujAS8hYhAPFkYxpRGYvdB
rgFl7Agq8Ti8FfZvoWNlp4/P1SJYzNtfHqyqONWV1MiMrtbRJewYHu9tKjrWCP3uIF2+6vRg8T4H
aKILAJrMbNy6IAMNI/xRHL1lC6T+ZgscwnGAFSaItki7u5OwnKTvBUHkz6zNs6yDntXcZ+mcs14Q
Egepyayp5C90iaukpBtR05VX19WG3MOuMtRrT78FfHi++JgqdmRI7oyPAyFvbDdARdbwVqB/DX8W
6yw0/UiXoni+XoBFMdCqSZtyOpLrH5Fno+hTqPu0VXVOBO+gvOQMulcP9enfnMGA+nmk7F59aqyH
qAicVgGKbmcNlKKzXQV1QJdPX6/Y95Co2rdFXcgrOstDwkF2Nj4wNrkAUHQuQEE2Q9HOZWC0TOO1
rZHZuGKU61o+4P4Jf0xPfa9wIIOG0zMc6hgOW/mWDspKAMRT3YF/biG4/LCjoUzjXmDbX0MV57bO
BEEEGNvzBJcFDGMhV5dH8MhWWl3v0ogoJbECp+5chzsnjFksnfLPh+RiMeG8QvWgGmhToeviQFWM
POIKH6+epqYD3OE+Iqp6QHVtKf1Xl35VwkccZBW6LzmabAXZzQhWmyMx4oZvHkEBY1VwIYYFGVb3
/2IjeHVtBNkQlkW9DOYF8xEzFvPjbXWBNuXgSK6TIqH8tvp//4z7wil2NRCM/byyqs5y+Ex2hfe6
AG6TZrIy1LRjGsR2FZjdhPfSSvfxOfM75TmU96xIG06CQloot4zrWz1gGMjK2kq/kE2J0q4Z5L0r
f0g0kvVaLGGLVoYZCGY8IDWNW6UkIglqkl00muUDcdfqe3HUsz6MKimTKdcjsMabJV9IKcRoHUcj
msBmnO8GigbrAG3JCnD0+mU3+7yKWGCNfdwWf1KxjMBwtwqeHwyHWmAgW+Du6m/Wg4bNHB7mM1ER
BLLH1DZ1X9xRe5zMSjWIcQPGHQM3jJnkwogJf7gk9Du6piKpXfKaRvALyiMUSVNno8nFRWfoQdX9
+Icw7xxhQ66NQNUMfwff2EwE1JmYsFeMbQwGMIF1Q5d9zkP510pN4hL0DoCKvMymURMCrxfY8Hc+
VoDu3B0RqDGZRYKhxGNx8Q8dla06QobF1irK9zmE8DCLed29yaO3qb2Kf3zI66fd3iMwJWg3vOBv
9MFdJCFsx+Tlj4N8LdB5OUIzAbCNQu8IyFOuv3t86eYcvx6CwP5xyIwCAwdX6EDPGYnojvpjEkkm
tTpjJxmfgjL+KSshFT+IdCLda6vABUAOKIteP6xjItqUD+74btLd/FkX7w8cLae846WXtK59pIYZ
Y00FwYpkbuUUH/vLUspjmqv4B68Xa5TtV/9Wx18NPWY5IHg3+RvThh9ssxoPvTrOntT9MSiNEuxI
Kc/vT+8hcIiipriJfAeAiVH6i6XcwLqoDwbHH9A0ATMclk6tvf14L41oIEmdjp4X+AeBB+ZxPtu2
nxzFhAfggmFnTazOAlJ9H/RksixWTding+0f3h5keW+cGat4tTKZ5WEFqDrQWhZTB3NsSh1chj0R
NDs38/uKutnhY+cHBzTlgp0YW4qB1suMmDq+z+aBRnn12belRviGGmEH8+RrcnpJWU/XhVjogaDq
TxNd58QohPltnal46NXUrcMRtOUWtZFdVyLU99w4Q5fboTUxC+haeg4JZoagsvHD/yn6lFUPA2rA
emn5OMOvxX7ZogVT1xoiStzfeVhtAB+gDYrXm5o6Rb/Ovw9mP6jgJ3LdCFfHHJjpn8af6gxuQwt9
PIJaORLW4FojB7wPM567Zu2t8hd/cI9RsUw48b0BUqEy502kGrX4x9YO6cBubuqdf7l0631vUQgP
YYteMQszjtfDkn32Rv4ba9pvbYqeXwNdF9uz2dHE2hnk3OPplVt1hmMumEb7ameqw8uPO7Se4gZM
0Wv+xD4zuTM5qfoerkre527AsECIY57iwHz9ufv9y+x4AWeoiEQESvU47IJFtsASvQVbDIwwln4O
XDh9gq5AyLuL6QNc3W/mdS7rzl9sPBpKNJG7HH5tZSMq7ce9pQNoibTi7/5R211qt6iHVQpYZiqO
WaDTwZC0j4L4fB0Wzyx+v7Z6cjAgNx/02WXuALY+vYQGuJuM9sM7499NNnwgsT8hFHAwCAkLtyIa
ZOmf5yjG6O6d4d+9uVP8+gnlRsGnNxIrxouQW4Jo5t/BlAJW+5/2qaGNXqkjUgJjMe4V272jGHxn
mLgUXLD72mfpKOtsJZzw7eKR7vjQbHrFVmiAxmeMUD5nhN9WFAlmhJXw0eNdvHj85HWyH7vbwcWx
ElRtbyTug+oGquUdYbMiS9ZoN8uoR39AuB1ijkWNRZF09Gc5t5wk0ulxIKUYjkTgu4sGKixvx4iC
DwdfDQ+Y3fCKoeYJVKLkoQQXeJy2xf3TAJ+PUSxpO6SjNiCPuSdiTYwzIYGgP49r7p1BBzM6vPRb
LU4dvO5QlOv47+IaKzLIk0V+yOf+JBd2E8FUDfVJjMgpH2Y+lnp2yA9tFHy01fYMC4pmvBqm1gpd
PS72SuR62y+UfJbRMkBk+UpGF2gvSuYxCisP69ISC9y+hIF0pV+8JvOpPsATKHJJttsQmYvrBUHF
gX6EzlkUUcEAVqiksXRss85XORSv0hGXBIA6MvN0sXKDFPP+HrEHzwll26y/Pjw7w6tlRHwGcaH5
yh5LcxIjNePntC5aHroH8XoPez3cSQAf6LW0o0LXTYeUjF18tdFtpu2UFp8I7i7wC3uPsT2Z8sus
ofppByB6h9jYvm4lt6Kgxu/L0JVzUqSkwoZsuH356yCLLxxkis6Eo3A7344KODmGAvbEcMBPlZD0
GD4wiiMF0l61H4hLyeyj3zrZgrp8sbeO0Fsu2MqbDwgzJYEzBS+VDHQDdewR+5NEFlCXYqZNT8YD
pvpLZvt2xS6q3wbFI1tpWeziNjvbn8Ry7YhFw8XsKwzujz/rAZFyHhozRZsedo3fNXnhwHjHW3FH
32PMOHhJr+bNmm3xgXsCG+usY/RkdHaMbAk0ithrDPPpCam8f0tF757CRGeu/eG7eSg7o+RyWFOl
wq9bIAkgRHIVFhKry5ygukCDpxn+HaovL2ESh5yK3TdMn6h6q3RI4ceAcNh21UYI6Ce2jDCWlZds
dVSa39kLfUJ9cBAV/4BzkXAOC30mlGVJfirq6gbim1K3+2b5uUOJjCw29AcBtE7TV0U0caRbSQNx
u11uyAa4McFfhwic2oeCb23bECzOY4z4LecdYAFFRhyoTV647sikM39VK+iGlnjvfbgJKD2N9xJJ
CMVZPIeINmAqZKfjExmYlKb4luH+9wOwQrJu9yfDeQJhJ5HZH5Kw4xzjHrIUcvEqy4DRMF9cSQ+4
7MWhRtw14T6gCyZhdRDvfEBZL+P64VR6kCTKW178phdot3A6BO3TEKXWPyRuzg3dUnfsrvWNrqGy
BuxYHmBoLGG8GkPjsAznYzEftz9CKvsXnT0r6rDxibzOipFVpdT/feq7t7cH5GRZ7J/TDs8A4Wca
lXV5a7fFUtxTR6N2/zaKBOq5sWjzfdQQ/UM+/ZI9IGIJU61IMER9qknBwzl3G6x9XIF7dxQmWyWm
QCKgVb0a0FzdOrvzGu7ogGemjD8jB07RHV2vxoK3OODtifF2it554eonmAQGKxv6PjKVFttTkpZ1
dhFvjfOARV7NmzTEFiiTZ4ZicxnaXLqboc5tZCufif2oBbOo/4I2k4RaLuZ3XSGU02KooSYamRDC
Ut7QGalQOjlXXnOBBX2dlokRNqUKUb6G+D2so1vyUYsbKJrLhQpqD3I/FdY556sV1zW6xfI30ftn
lA/q0oruze8doGFqOjNc4edXx5pLEZJvtAsCjqCFR5UNQNBmpzJXkcEWWPgc49cUDBorbkcv0bWS
2UeQsFOJztQMta3Jff+eGkuUdZIjoaWGlrz2CDwmQdYd3DL6f41Pqvsm7Ku4KeUeKUMrZTK4TSIh
+tGctEOrg3XwZWhMFkUSjLSHuYGxic5Af6qcXasrNejtpMUE/iJsiwWGBlQ0xA5YN28VT9qnfRBe
tNAobRgn6ZoaYYCLGQ32E/UJQPT9KQ/Z8jXXUj/hyaGjE+3pxGK+yA1i5sXDjbtH3n3rmnhm6xPv
rWquKNxQ81EzKY6Gm3opdhS53QqU5tvVhxX56BYWy4VcR99b181+0U1BWd4sBtXE2EoQrtubSNGo
jpcRxGWWEuFpDK2TRjhyuWy7D3tqxK3e8qFfS7BuGkhXjhT0kcWqIflPTUosCdDZ1FMT6YvvFdtg
lCd6cTMlgk3RXEm6OqB1yyVhpGwNKuwTVFjMkZBI0YIDpHw2cPjDSkC6QAl+ihlMJCnMIZR+XzE+
fdPzOK4ilyMM6x3B5tSjaRl6z/IJ0V7OGdK23Zeeke0kysfoxmJKPvuUrweXySszlVLz0SbsslBe
Dk8ZV/vav2OsOBqoFwsQT3xCZvigaJHr7jJErLTSnis+SIU9RFkp8+k9A+47duxIzozyRaVYRqeX
FKUmN5rLMPPIm46QFEiYTNPOuRmZoqUhHgu6wTdpJ2uyE5f/LXSdfGAqpYiEw41/B9ZqcVFqbce1
QWx67BufHnoQ63kPeBzitESfBgc8xWWAu1U37mHKVvCXQMq76mMboSbP3iZSHXgBHCVpun/RbIw+
AsS0htmNevF1OqvJKoN4FaLjqfXZ9A/1hYqV9EqgnmVqxVdM+yrRYCzoZVMSiD94LLBA7ZEh57B8
x+SuwKosrK0apot7x8VX6+DZlDu0jAap395D2w1L3L/eptSXse06FpZ7rLM6ypMewRq1rJc6u1Qv
AkH838BWCYGVupWCa9MzihMdvREZd+21wJPVJMFJo5Ouiba+9hJTtgAkJS/4boWcRS1K1D9BSOZW
p4w3TkkHQJ6vaIMlN0UstVTmjUAo3KBQBdRCgLzNISQ/jZQMt0UuqDwD2msyT/ybsUpJXMEh0GeK
bil/UsdOY1r/cyuucaMSyRJuULj8uhmdpqWfub/bZhTB2h53NM97FRP5IMy/IiZ5LN4toVOq/UQW
8TdX4xL9cVySKFafjq6gVPTwu33VK8tnW+9Ji+wzXGFHCQFoHDMIAY3tbj424Qybym2h9I29q7pa
lm3YfonuaC1mcB7pJFfbeQexKHaU2qFvpUtFdaAxUO+8c4tAfv1vluartm4pf+cwk1Hv+xqx2Q0D
o18pXbA+g7+zqsxcgqaFg7zHsxtBK+QulzWRoI8hbpQQL+/5kuJvuJ/cpa96eOTm2AIobpHrjXem
So+QeFsww+g+c4TJMbRowuxbDjultQ8GUKwAjcCtbxsXI+jidmy7TcAjJIIiphbmZkLMMQSAmz0C
PEb1idJwZVJUcrTZXnzS6PhdU5YuBtCyB1xU4H1U96MrYn4U13xE/gDXNHWQ9GLgdfwfQuG00Mbp
fN/U0/0Gm7amUDIrpI/X+jRSfabG3j+/RX+u9EikQ7lkBV5DKixOCmbzsdnUbVJOU9AuByOfTs/a
T7MvUuD3e5ddgvY+xWn/exIX7NnV3n+Vb7BUXZFPtFnNsOqTEp3ss/gq8OvXT3fRAtPKQuV415ct
gktZIyS3ntLBF6A37LTfdrWr3TlDw0zcCtEpN1e/vbjQ5I1+0pWFoJ5NGRhLLAP8gsttMFs5AnzV
QCNJe/DPbh/URtgbU19UfWzepfBML1JAMktYLqA/cwxxMtSOqQftYXMw/52IpuwYgXYR/rxitaAb
4qiFryOSLqDmL5IoGnQaMHfu+6HRQ3CyRtMArlfy18gFe/vOHPMglluUAe+8KYEtn4RasJ/HYevi
izyMIIUe1MOFQMsk828/0vxBwpf5JY087H9BcYcJRmwmggGgSKlgoZqnK2S8JHWls/dTUqIqKM8J
a22HT8RJCBc7zdgue3s3LQfU2JmWqtSVcdL4XND6a/Aic0WjO8RKiVUQ+1ezmP8rN+liDRB5ANpe
lSJ8SUZC/Vq14wGJobU7ROOKgk7qS8I3yVOy9v+BI+vWf0KGZpBCL+5ziYtDTsf7PjpZ2u0Efrzm
84Y00FP0hd6/GCThum0i0ZIMjZTzJvkG/FkJqsi/ohxVHAgCFlYNwK2cO0b3QzvTCS9Zn0WhrOds
bLWaSHZRm8L1TFmm+Jz1hVKSjpDeivaSp4M+/wDU1n90YOC8BU82eKlFpNp0caAyAZSCgwFcpVPP
7YQRTlj5oP8TSrSqIGKEwd5U1DKY3XDJfMJ5HY6g2EO0wtxlhxASoRlGQL96tfkfBBt1d6KHqsGv
tj8SO+zqasJ0hSck1dZUZHpWZO3ZJEOfIr5uUFRlz9OOBIwh8kY80tVSM2ahRfTheajJ1ZqpW4x3
VWoLWZhc6OAGCKmt3LmAaW0qu8KAczdYc2o2bMDZ/UeVqxSO9J8HBx3UmzWnJzinwdggKxwq2xY3
GJ7gPWRCz5gfOD5BvgSgFitU5xeY1IxFvTf/jG4HKk80fWs+lVag84kfzT6CdcjVXZ7G5Rjtn2kt
DxnuuLWQvN3iRCm7J/Z2axbpdYoMz2Hx43adXVkuYiiu5KDt0UbRgXTaoKQtt3maRfKD0phE7Luq
+RGnXWVrCmjJ+RaEyoVtD07jSWPkvTnkj1sBZl6LQYeNbWMI3jGQBt1ZmgK64hUnkwcSTZ21sy/l
SFNdhL2KH/kf3rk1OzroR2wKucC9U8vhhhpvVTNiMF7b3M7142UuGP0KkY1DHtk/0oIEx9vBSc/K
WuxhZCjZBMuWr5h0GZFSzIWgKPmnFIkcc/d2AOvVwFDfT2l+FPx/BUncBzRJOvPReb/s7ITbbV1r
DTsPN85qUrDUO6rPKDWWdqCC8VeNTop6g4SAUo5npV597+a/enbly2lUZq3V5tG17vCDn3veZUE2
SFqKxSsVJQ3E+xdlNlyN7G+F+uEnlidnqpSZpv08uIQZKJeSZ+emyyWMi83Td4XDNbEC6juRXDGM
2oNRO1tvSPzXUhGVPaHiCgivkfxs0g5EPYC1fIHhrOkCR/js9hq4Po63VH9Fzcprx8K4/xxeY8JB
JoiOCKlm8ibtt75aJ4DvEPG6R4fV/GiPBfSrhqcP8S1UhEt5dTKASxY/CLas/d58tvGG4QYiemqR
irHkL/WjADq6ZihujyS5s9608Xakqsh3Bxt4E7CYrH002lSNlUj0fVRfQwAskXhq8a/qdpA1ulQi
qMVMEAVJIf5mzrh2/luewybgDA6YxUIah12+BhSJc3/bv/F+pH8p49//hwe3ftKtgBxrjV9eWhTj
D8xAocRmgs6r92RWxpQnls+CO+TY3HS/IjsdeLhkzb8Y2M3rhgpRXaHweox3KJVI3aCrgK5MGCmg
p/UTVyk+MAouIf05CKoaE3Q2O6GuhHY8lq5vvUN7UanSvL4XqqgyUkUPeQGEc1rpVMGPnY7INUL6
RFGsmXci0F67MNpyCfZBL0De+bonaOSiltLo+epGCij1QIYxVjdf9vDvUtZqRaRCv1/IDU/AlZ4g
tLWWS6TyC13DFwMvsqjPM3frMcKXToam4ljQGFY8NEvNt1awPKx5NTSgmbzMRvRi7rqQ/+jwLUeK
3F31B/4othN/+GujVVYFeHJJMJFozWZ1stT/H+RIAYSC4hON1Hxr2igIWYBz+S547HArUuD+fAez
sv+xiWJx2xugES0FY7q9Hi79JLpz7tqcIrpKiyV04taiUEfiTY0QEqShZrzKJiQsfjY7P4FBwyd0
JzlDEnt/GWK2m687RbXgCk1wZ4/8H0bffmbKrSAyvMdHrCzEHjR6plF7sRBTGJXaz+s3JTkutcrk
OnWLLYeLmPzEXBx7zQFtcQ0siGVnNFyKPswMWcC8tNz2c7NcUzubNFUwBpFhZqPyoZywmKhoxKIi
EEJLm33Sysbpf1r5eRihjuHJnFBt1N2XzXNGDhW5jghyYKedUdUiUbPXzUbWC+RcN9IBRpCa5Ak7
lJb6mWE92ragU/aHqcRymRTpcFRdSw1HhuwmxXmrw2D/nKgHUnRBbr9g8wY+7zWFZZbz9lawFJtc
b3yc3KyCEggDiIbRsh1YOIypJG3nRkdlobUZCCVvWlbuZ11OuiXeBt6zjLP6Ko2iUBkZ1zWAGOm1
umYyHPmSGkOmliPqUCs1YAYAmDssvx4TaK+589QveiIwFK8VKe4qcWYUViFqd6dmfk6ziLvxMqUT
d5bxA0JHjCtY/snlXw4EoWVO7M99Hhy0UAWHTA4/qsD0lKxFsVrLlykvSWM2/BkJU2HtgwgH/qug
MoQHFf6bKiKwMgsTVp1FCJaLtJKaCSXaK+UMy/TVbH8OBcTJgeDDNZySH1mnIw8zXf6QbB5aX5RP
m3icF61GMKxMQDaHkV5MJ7jVO+Y1D/SZbJDM/X+qIb/bIs4m04BUFTviE085Q4jNpGRykyoYfm/u
74BbFaTevYAQLnbDEczRnx6TUY0vfskuv88LJW3FR/5BF5cyTsIsotF73gfY6hsVCCmdGiPZAvIk
3OJUw7JdmBB0H/TY2Nb0JKNU85sHvdBwCzNDp0JB1m94R+gpiVEXqbrSJns78qg31+xN2KSrlk9O
OaPDTMGVX7uLylVjdizxHsTmVRWru92TVCmuLv94+afR1EtzcOJwb4u8ESkmOHFFQYJD8uFg4v+t
fWkgybVXCNn3Q2XHoVUyTQPnNbktNGAtbvpiswDLqElPlnKgMdVsWhvSMG7mkJzwaN9BRcFbTxUr
Fwy1kJXan/NzEZ0Se5LDZAGCihy54G1LKA6N9kl8TmzfgDuLoPn9gV7pNg+TDYwC2KPtYKuGXta4
dH4WFJPpak/w/3hzENxFDojU/VmVGuCyrACYOdEQnunBdpxMkvTw9bkZUVunXG5Gb+1srr12ce6D
GxQZyt0wyX5Vy9eLGnoYv5j6Tu16fltzjKJQuYGIVtsqhzKR+U0oL+UiqclYfw/DPUQ3Trz6AaaY
CMZoclgH8DRUKW6ld+BCyLb7QUtm8VgGqOUjUhampg6+XsMUd5NFa44jgV8b8+2+tRstOPu8aNA4
E8Qa+E/ZieoxJRmBQ4+lYvR2OCrjKjiliwkq2PKVf2hrQtQ46nWC4L1BAQFdM23e6UvLHosnRZti
KcnTScWFCQSHKZZxnTKJxP9a4oG3DbAdK63zx/GflpYRGg2qm2HNJPABlnfFYpakGEzKdvuUXqrn
XlfkKEoTUVWgLj7hZelm/wzWuk83V8c8Ayw0XRiWnWyplKJb2Ra3J8n2CWDtdGhrwHgrMnh7nDXX
/PqR56mb5iGnpS5OkQc0gxQw0Ree+nzQddAzz/617WXy5AAoSvQy2SP0pg2evWeYBsqRfEQvahFz
GnOlZF8ChvHA3QJdV9QircnuO2CSRvmw9N4gqOPZelC0fzrfkWwaJPTMwCuI6c/U5vicFaXng+WR
UXrFohXi1vZ9YNjW3WtrUVAUzOKHMftbaYMb5CF20NoTXO3b63ReWTXCqSISnImi5ad8777VKdtG
Lqgo5QMZbB4vE0r87d7VN9xfQGF3vHP854tJ93IhVowroXoqDYtYMXAV9+sXebfRkOTrmyTF96dh
ui3X/DhGqpHvqg5xYaxqrYQdquUdtCChZd7d+rga/KMSVuV9PbGZ1ZejUnqtT+xmhGwr8KPyGzvS
32Wxw5aalZR/PXokB3sNHYDUhFHeTovGnUPa5f74wDcIXriCEyAD93wrRjV+5yAvICHTcCC2a/tf
RjIroJjDOZhclgvUA6l7FrUFS1I968jSyNIZAFlp4P9Niz8vRK15bQJ/E9vn8mRGvmKjHgPDlU0q
zSF3Ld9BMzFl0LbCO3ChwqHQJ6gtRQMLyeHmEgewnTrhEkWXMwWc7qGF/N8t0d+i6VjJ8GpToe0g
btIOEHSL0Zw4OC7WJm1jdZhLxoSJBdfpKG+2+zZZMWqEbSE4d9ycklo28LLgJckvxHVrKQZhAHJa
HuZecg/yvYQ2f+MfPWCZMX9nwwOs3sI0FfZGMeuRqwVaDWidRQE7BftpH65JvZMiUBMiKDoeEJDi
CcSsh5PPs5D5uM1aBz4pkXyppjlSWib6yeNDN7rCnk2bHyBRe9AmmE245Jc85nl0naRBN2IQvO5I
q+NmWUH5MW/9+oo6POf652kyR5eonzoXcuxXm59E3zVMA3ARoW7Yn7uyz7Moh98RuiH8pJVZgM8m
xxaAKPAqPGken4Vz2LONAVOnfg+fGi8hfxWQml0Y3tmMjU/Y+hYdCnPJ678lBcq3xLGOKE0+bVa1
FP52zifgIJae2cpSy98FZQVMeufWEUw04AhRsTB92R8a+JrxcpLRwujOCJssVR0fBKWHQ23agufD
N95MxGbyvC1PWwADtMpug2L9Ai+Tf/YMikJW3VfDHIa6WYEXpfLlQAQvrKrGoUFr1o/z3cQbghOH
cmha+bx/LJaMxXyOklqSFLK16b+JS1NdMvtc1Zh1zFv31i5L0DvE+xhE77WkBSLFYw23t1O3kOEQ
YhMIcnx2XJHIOk+QEE0Tp674pr0wWwFZF5EE8bZqWtOLub+JXwb7y/Pz8JGUIu+Eis519SKw5hY7
wqs5cjOepLb0h6l/L/5VcRaXVnPT6JnpHYIet0HHoiaUnkZuQsN2JKwMwx0SO8NNwa0C9elDh7Ea
hhoKQMwxXhf5uCCfABhHSV09PFujwZ6CRy/2eXuZkZrg0QwRJWB22iu//8yS/sQX5Hn7VcEfraxG
GP8Y/Fiutl6CvKq/toPMdvx8uSBl9zZaE3GaOXPBKa63Om3Z37hWA5QCkoKHVi/twJjYvo+hSaqn
IEu9Dp/dDo+5oK1ZTrmVIFcyFBB2w8oa6Px9hUhkwArUP+5K0VeM3s3vr0RHgMdTBS0V+Ys4cvFk
qJG6klwK96uGgIsEzgc/fhoIXvP/jIcWy1AnuES3wDKJE0XE3xeuK++iRK85GPBBBF/6aNPs9mHm
caL1JMzTThIm2vlvFyAgh3WktFUKet2MDtFqri1w05rDtBvcrtcvq9EuRyCUxSvX5GPqGiFJIiwI
QXMa/pHBjAtDDx1T3UnW2XvWhhtYP8MNpykBHF1ZyStn2D5Y3uTcxuZpKhith5vUl7nLDNFGDjvY
891XinR1tFPf2fg8/Ickq3UgP9Yyx2aSVA6ZkTTeF6Ue2Q5dWPRH5Kk1vH6cf/KUpRoMxbfpobjR
CnkOry8gMroUoyrnEVVAUxGR27dd7CMqBXIabQ9XaaZvB3/3LQF7NViUEbdfKd8ZJjhczWUeuXsr
y47f+/ctKo3IejgFz62fEXJ9zJqnkIVe3NVxJoQWGDJajl/5IPmj3aRPqw2Aw61TefBmjq3usPLV
7synjFd6WLWN+Q0YGCQH0NYT+cRnp8WTouhvn7/+RsVI0WPrIirPHseMssfxT61TVuPbh0xtNAgO
2Np1h2+3vt1pUAkvFJNZt2azObmTHcSRjWy+l5ApXDfkQPNoXqTZCW6xEVYiKBS7T/BemNK+mvIj
+yJuyIEqGPDsFQEp5B0QA5VDpdKkFkKzB15SArGmM7vAMxmQpcquYVlmpf7Ju/MRpC8W/3EexedE
3vs6emgpKrBEnIb67E/zRaQCdzZFmaaB7aJYNlgYzHGmmY7nG2W/bi6ionBJVENqq3ka6TPsdeHY
UpJobVbmpG7maM9V9qEL60F4HffBw+RQzrIPzqn354mQDXGuxYaBwzYIBuZOjBK/EubRF1AoxJ0e
NuUTsKZnffxAVhH2CBZCHAsOA7uLobllpWffep4kgtb44Ihc1az9u7FINfQMKRWEgcKZ3LnZtVRi
aidjxieeJhUveHN4bqtfSgzCcnsSRqSkABttozywiOGv3Y1FRxnprbzx/Z1nA+fMRmUKWoe0nihv
sZ7/vnogBP8tKJU+1KlC+/qjRCOXfWJpAjE/YhYBoWUEiir5OpMCQXfbmmGW6E5eLlSG6pyRr7v/
Uo2vdAtZnIg97/VmvmlSOsPHHRcXCSLdgnLSOlncq++h9dVaaM6dZRlOkDJXKmj5cl9R9gQ5sfpU
jPk4KvsrsFexOIW4USIIzMIrpU2klpb2kQojtpaTcNli9IbipmZD2XrxxCPMeS0dITvQShvP5GHN
Iecy8AluF9KzSg1LhkKr5DOGXTiTf/7x0gqpF7TXQKQUVIkr/SbkZIv++qgAoeCt8lpuE6/1coLe
1KP5iNyDBoLiil/CHJbf9y0YpYibs0If+qNgWo0i/SoBsy0wp4WB8oS3VhWhMRAOt7fKQKozap/M
80mF5YgeCPzlRVZLzCENL/W8zx1fxGI/i1IaJ3qvibMXcne5Wct0SpO7E0HF7xtoVAhQJgQPiyce
0KCCgRc8GneyDzLYZjdTdkyZi4ZDLRQ8ABHBS3cqQawCdiLzPmpevc0teedxztkrkNH52iCqWAmT
nsDIlR1rub0fVytJ5qxduOPfOwAeTTXzKySv/dHLuQyqelimeKb6wDh1NtEb5JksISNJv1vO7mfF
MZXd7nj//WfnXYKffCdSy/YVvfFQME86An3xmEh31kyO9xb3XoFXDxy5XPSXPldnTo2RM6opRW8y
0bbZ1GKgqqD3vL6ZQYNXeBu3oWoTMV6hxZPepAzkwwuxmDVwRTp2i/AKhW+wnzt9Y/3/+w2NLc4L
3FghyqAnOQe/SNKflyDZ1CcsPMklnXQ6aedTMMiPiJqiLFwKCfnTy4eWkDozJQZgbY1sxXS8OZMc
s6Y8uq9u3tfgNCZKp91+ZvdVCkBn7Kv3lCbOQDzlTp2tc3V1kZOsMGWX8HKlbYE1V02kGDBCxv2y
mI4youRgPY2bpxBwFlTR1jKsI5Qbj+tj4cogaz/WbXb3A7Dk1+MCztYyCv4WWkHwDs4VSCX2X8hj
LTyFLtQuK8o/VdQkXhauwQQqYgYIr8MKIjeb+cyJCgJMMW09r22L4AkSI13PY/Rnrel8YQmpKxZ2
RGpPlwqZNfk29RBewyVz6GDMALdf8kwB5k1Qrngln0RypYe3YHEJrndEUWgfLq7J60sQRZf9MfxD
ZYIGo4VBa3R+5N8Os6vsagGKIJRiXVjxVHbBysOUCQlZy6dZqZrLb3MlGGtPj2tJbVPjF6hx2CGr
FTaNNjpPg0vnMaHHAxFkfclJ2n2r+x+q1hWHZUlDdcqLMkjiAR50E3H/6s9EgjZvaONsV2YU58sp
0IKXSTAfACdgA4omkFCv5Fy98tbkAMW8LFFqJv3kDEvtaBiXKslDTf9bKzeRlzjoKxBQPzd5cYLy
CT0wmOO4KM5yIvG/+ODl2hQTQEdOrMbseOvxrVZ3bAn5U5s3PmvgIGRyKWqWPxv7I6IO1lkkRaQ/
5DQCGOINmJVEXmjjs2Da9/s8bg0kPaJrnDTJSUtXgluL8ZEKOHoQq1CKHPLyjfO+qXsaxN1xHOlb
eryuoYn3AmxKAw8MOc/dqWet/IiU+kwIzXIK7p8MEaULiGdxqF+G3i1zk0D8wkGFh+s9ahtkTieo
ZDX8QK4P6/yzPe+oEgGnSiujDl7P8oGC2rqWovx1A7st4Keo4cznacKSJUnJPA2MfJpmKLuDmNcn
dqjLr8v8AUBg9MA0DXCFzMp3ZurYPXp1VSCs1oZx5JkoxgnrBi/PLiS+Z4a4V70LW5PblkpzFxd8
Rq9bEJTLSp7hYwlxnKuPwTnpgK+cjyNRROrD0KiOm+6DKwQdtFnB5UNwVZpKGIHKRU5ddEOygmPw
vUlDOJ1hI3rQoqDoGA80X85xT7xPOxw72CiKIMPD4vj5fjj2Lrm4kuRpvm4pLUMofSD8r7vLsd/f
GRGofr3F7Vbrik+FdbZy73jZqK3HKJpKgMPTn/eDg4X5kcXCMTB60bL9b9r2VFikOSwfPgkpA93q
hY5CQ2D/f2H7RgprM8DLgez+3oDtwIuhumHlSRYQ4wZzTLxiBk8OlK8CDQY4ZtQxH5Rmbh4nqTTq
8bm/ROzdE8FOzVbWJrxIXdVRBcwCM35wyaTDOFJ8pp6WP4X8kWkCfS2K0bY+U/YLZZT4SvML94tG
t7thCXcOcZM68uVA4LUiqDuY9+T1LbuKbgihqgZBfLnes2/lMgRa4dwwphlfqrFh1lFycnnuNBT2
5Qp5Ke4MT53nT4jIJePK5tdacbycQybt2mIyinHVRj7l6DJkawGIQAEnoiG4tQX45bYvBgsaOwFK
fd69KW0UnFJGPSUgTFOd2/BEqHOxOLF9/BGiqwltm1YWIpWmj0uxiO35iLLBmfvm1A1LVijoPuOo
Ok44RwQyUgCieKROof85rrfHthJWUq0Qct3rzUL6aAILEAt14L9iI2wCMBISl5qyqFMjchcVD9yW
YLNF8oSjkKHkDG+HWkXC+k4NjVJDthsGVB2djufuzS5atAamzNSVS28s4PzAfl1FiqcO8re1nb7r
57I8JgQ+jmisXZS1z8RN9TW4H7limH/L7ChKQVLsUQwZhaFDkWDBLpnqxjVYT6xX+8IjGFh0TKpV
h3RK9JUiMD8nCI1RRq/4AagJosMo99aJ1vl40W6cSTHfyFBOKZ9XwcbO47FUc3qyHDvWhkL8pOcu
vzPTe0rqCggr6QKLHm9NJp6hZL2ePGir+FCXt63sACYzzTIK9KN2hngwJLmVtJcb38ynSOTepoB4
HAFIKCvezS0nIf5+dmJRC1NFvZ6vnzK5mHcgneVcURAsaacy4Qta3gopC8RQDSwcV9gO9M7Luyu8
KIzujCwKVini9HSgEgkN5XmdhZOzo+opEdIJqpHPD44ZAAYxtg3nF2FxX/Ms0jRwDOQBKe3RCmim
kw53wwBaQAg8qbsnc4jDtRuqW/hJCABHxywCki/+qpzld06z3Hd1yTVigUN2Q/NnTfg+JVvQxRBz
2vQOUHz/bzFqEcSDvOPnYYJec6F1XCz0446IbBLA+dwIHiKh+csB+DwL667LJsvRocdby6Rgc93G
7gNSMsjMwMQEIm7hzvyMrtBkxImI9bU2mMjmKYCz53pvm2ngPAloy85T2pvZp3jmYuwG1gA7+pP9
J3KAqBjO+x3br1WdXnfWooDc96tarhzE0Mh0WvSt0vwKmmbcI/TFM7o7BvOXuCysyGZoQuweqB70
kmkvbIzTwsvHlXOR1uacRVa8b8l5ws3OSsVqJ607yFpZMfq1Rgg6leZf2ADhHGb61vtZq/9JgqMv
oy89y/32O0jfYl53b3/kBjaf6/pGssXCTMC+Lm+mg0A/+mChQV6jB1dCH/rUIUWC60TxkvVOLYi+
rqSUZYU+T+yRZgSgqmZCXfG/RuPWLaNXPS4CV+BVQ0+YhNV0CBVjvioSkewJa56upzK5VsEUfvD7
XaHB7m6mFygKM96+fplARi+zR1Tc2EqQK2fltVIW0Vn4roBw/s3ya/HGuCu2NccO9SSj32CjT+4Y
iwTBWBJc6YsDibQw5TIj0Jk7TnYKbFmyUCO2DcBvRUjYcRc2jkWWF6exENOqFAQ7A+/34w8Qcc1m
eHeJXcvaDdaeDxIZe8N+ecDZ8vxJTdlXKf0VO1VsgE/lHIw/x3Svh0aeF9PAJ/kVMhbL3YW0d8/J
8ndXNVG2MSTBFKu2LB1Bm2UPcZIbWSqOuQxUZNCNidBLX9G1h5gdlWVbZE9WBLWwLY1YDg6Qp3iZ
AOBneedqVGZtQoC5hvSIL8hOkZWDdfyAAJgOenlwBgG/XlWg1S0b1AFjZ2F96/ZgcgO5LYod0Nlu
zZiO4RaqAmYxxN4jRwKXBqzMJc9/w9ovPIyi/PNfl7BTjfSodtiy9JIou+1jlmegLZpv4onFYJeT
m5sYGVZxJamfC05H/RBaTogUE9CkeCEkxHiZgEMzML/3Qaa5+E4P9HF3BJ0udbb9bL5d3R5N6QQZ
jxud+gIR/khCj/pfbzq5UQq0biHC4GRnh9p5ixxpN+eDUjY+6RiIcv2a+4aSJwseUUd+b47vp2r6
zZPqpUJ0eCCAlW8MDEhSYuZwSjx7P5hkCnjqUnlmbuPKxEovkoFZQSGncytfPfXUGQ3TpmnbECUq
bX4kJRCtp2Fazew9qtRMZha4SAFOYRF3vw8TYbEt4HWgdwbyzYoXnydUYK/9ifw7d8lq4MpPNnxl
3YXiCsXBb65rs6ULIovpWR4NusXBNoPG96BAXGeeYbc0O8h8wZrkKFJHzrCVthpAYkvO5e0gEmHU
N1YfWw3pAsZqF0dFe44UsRCTdrZeJNLh/EYm/q015yRAlO01tE7vkavbX6QzqEhFxVtCp49uBEtN
pqhV6GuFP7Je6FJgVDdQ3tSjk/ZYqO6sdGmQgrrKXDE6DdBgT+nrWzSdxDSl5GpUs44GQGb7NxXR
zl39RUrvc16uize97rbgFmAXUmgmIXvaleS+eXQ7oBaOLRzovGkEAMND/tlhWv93jISfKzy9RoQH
BuxGpaRjfWpKt6wjWGjDconoKH20NE3SJiTIyMe5I0GSm+R6IjO9ImDth5DAo088z2RDd5gc9KzY
Gl888yo1x8UThgNHW5FwF3jNJ58uIvzoHW0e5PDb1ky/Qei/79JsBoFAzj0egc2xLOCTI5QaIzYn
frAVbnCEqMGvP8f4osw2wsYCjk4VgWzg3OyEPx4uFQLkfpNGlElsW9eN2zX+ZZ2crzbtad22Z9II
pYkeW/lHcPYoVeYEYHXPGlzH+jfFEg9mfKZ2LwarwNyMjwdEJtYiRpOFdSiHjrKcpzinIM9Nk0eG
6ejbQQaJAL2I6dPkbZdy+pQJYzaEKtEXw60pq+DSVP+rXjtYHCeyJNaDN8o4Jpf7ECYUHN4I3LLo
BDh6gOcGsg+sw0zNw+xZ8JKSPZgeDYov3FqlBD2sGpJ5f7aOKCmeXbNUKq8PWzSO99XKWkdyPU4/
+cttyE5+nojGA5vL5RO79qQ/9uOFViEpQPe8lS/j71hmPg5lA3uyfQeb+V30ZU2GQRzvjbA5hvxh
NphAiSB3p6rPP53HIHzkM/V3iXYHvHMt2N3IWGhLGaT5LRcQdUNVIHiQQlrTrN07uHYIguyF9BR+
bULy4/UJNA+BlNLorKb3Ux10eCBEstV/mZ1OwJlnt5YynDSDNF2ecDxlixGVAmkBtQb47bppZD6h
rpsloX3S50xtxP8sF/W8fCQBwCiQ+zz3U0s3b9jxakMWlqPMFef1ApmSx9NMWHKC4WDfDpYsOJjc
YMUXDoHBZ6F5YstGeD//0mD1A74rzYTEDBUp7OeJdXuaIx5JnWGWkCDB3VkQrzWkj51Rn7mxOPxm
w38evXsUutBAHG5uubM4dlADzcmvfS/DJZ5U7K37b4fGIO1Sz+wkOvHSMd1+2WsDzEoeuJ5Yv652
N1QY37Sw0rBzjPAxH3/CEIV0jngFw9TPQt0n48+I8qC8aDl/Vvr5d82Tf+JtuZTQ8gdZc7UXqUns
yg14I7dip61FEkh9SKBC3iRrNbn8FGWMWWRJDSGBad2FlwQCJme8DH1Sz9h4lWVxl7AWl4KC45Go
1stoeBYybULqSO/We37ak2xbXnKQN/ZKc9Y0lTcpMYHApmcW9N8php/Yt3f5UTep18S05NvOUZuh
SE8+t5wMnqhBknviRrcrrQz/koPTebcQ/+zsa4r35E6oj7Gs6i1tbCsxppbfbYIZ3Jnloa5m7Lmw
1+kV+uUMQrhKqgUcjL5E1S5N/bETHzyYd2Edyg4seudFYJr3Z1fxpYQwhX6C94WcJ44bF702CL14
B+dNWMBz92ZZiMttnVcnQbdo16nePhzjYPNTT9yFwmTm1lxQCgILq4DpOLP55Ie6sYKh5BcS7fGV
d8ptFy7uqIqk3GUlBi+Zwi3eNnwKyTDPU1OhZyVldBZfqLYrGn31PVrXTfnGeS0iOGj8osessvZJ
gXpMbqgL+rcOLUY+TNVvnp+MszUONzKn+vUkvRmNFWrY8rLgvtnPgpUAq5dQXjqklygeXfRN7Pdz
8RIbZC3ac4kbcYRhLaHfaTUXXDcCPV9J0nujiHViNrZIrhJUpq0SJFjtwg62WownnTu5/Jye0JDN
YyxGQ9KoPPgJQ7wUEIHocaY3Dj7PjlvgDworG3q1zJhxtt9481FJo6clCAynVH+G4VwvS+yKzGxo
g2fGN6kGNjxOIdlIQntmgDHyjbUGHfCIJs+tIX3fryNc8Xh/UCwhqmaPNZud9eeksU7rAZ9FovCE
Z6m1I1XLPLtVPlXJPNJmHvsdR/yLDmBnT1Ug3WrubtnLKyEK4JggMn9+/ABbKOWhft37g3cBy5Za
FoA7w5evaypUtQfoWV2fZaYiXvfKXv1mE5fVr/11G91X4DR6xBA78uBEbszXZexp3fQOjm0WcqNx
1rwjx443WR0kVSLqNeq0uhuItkl0KMnxYhnpOavA4aIDdXUZzuBO3YgviIHJi1DEq13lplYI7M9/
adaaRPBitgMkK04KkKMlypVkIMIQ6RK9TC4HEMTeuQ23CvUZ3FSUpXjUdsDA9OwnDfOvmsgdoXy+
7rMuncgtPeQixNKZHwcT3CLfQcWGgwGnDrToix3WPBUg2/gOlabBUIMa13hg3wIEUTch+pvAVmSS
m8B/puexg/mWe6/qxMnMl7AYDTnTeyDUoFkthmkDFx0Q3e87UGItRxFN3CFd+v7tClkH//Tf3fol
ncRLuCbBN57QVdRniA3vFbCOz1pT3mnA8fJovcaQcBsr4GaNxGCbyiPEllXdRqyrwrLHR/7OGkBD
08Qdi7tEBnByHabSQT79kE/SLlUG0y/DtV8foSJjy+bTVNCfeVPr4f9BTb7mpR5AsKBSN6ippCgC
fCoAD9N9Te9arF3r5Ij4Fx/Zc26nvGKMzB3beG9MEvJ1WaAIMoarR+EAgpfN7DDyMwdZKBKGBSeP
7rct/z8Ugh6Cp49bX45LX2fhU3Pf6E+WxL0UjSQOmfsjJ1GYr3f9111WN7roZAdeOABGH9EvaKWv
a91iXGFUOQBlVUtJgfhxlLf8k6ckGb6BHraRdDC085EJOBSM8IO1ix/EuRhlMUzt1ivDuxlIuEK4
34g6QU/eZsNT/PPpxD4i9M0xnjNvMHfUtlCxLdy+HXYp2RbrmLlLXNGVIBYzcJCO1S5cimkXb4K+
0vGTL4q2/J6fVQh15l1vAqHMQOWmWgF+1etohHS5NmbtpDAiiIdq/OssGjX18AUKbRw+wk7pSNW8
KAY3hmcHaG9/pqI0+oid/66SFSj1EwJvy4i7DUQylokd14Fopa7VW4D27YwS+m3k7I6wHDe8zPLV
ZRic3jz/H0x544uk0PL1T6PF1PY6In4bHYnphuDkTWjGvTsFQ90r0vkvt1FC2WO0e1CgV/sk+q2V
7IP0El4k+uRqQRX88Xg66IyUBVml+BSdQpDBuPwaTvxu2YhbGwEe8XVcZ9U6G7lqtMwDTpcfLyl2
iL5+5ZP5eexgC5MAJX1Uhp1YDJeTUIXsGPDNq7xUH+c/f/fxrD98CXy5YJm+PuabkSAv5yP7V/qW
Uzf2mDj8cRsIpgoy3t13ULdaeZD3cSJ1QG1jFMHE28NcVn+vaR4DP0n/PquR7KEh0KtB9NuHfFtN
5bPm/F+IdruNLVdKwNwUKGsIcnmI7siA8bKd1fMcxp8wCWLc5XJy1XVFdHMTx39WB7+P92Cp9h72
d9YBmZJ+eqVrOUh74FlnQT5BZECjFey3ZYEDcIVC6Satovna2mTAbXQk2QJLl7qz/4IS0Abizl6L
uQFqGozUfTP8/Alrjn2Ved3DSbBHGDEjlV/RnWfZemiytDefxnDpnBjynxSKH2k5m6nv9Ob6mBp9
EXtztMWSP9GQajUyRWGbxf5/3g1NnQbvUquUfen9LdvfCN+jPT8AHqnixdvpXC1B8SPyiRfasSJO
+8GAu4jCWTab2KODn3ybI4hphf5UAVtLBwHRD7HHKaR8ForQhDwu2oI7u9KLDA7ixoDz3AO2vwjP
kjkHRmOS84rm9TfTMVgDmDDlQII0oSp4prxsi9Pk0pUYvvgUCXvkL72AjPO03T44w5vkpYtZYroh
29FX5IXjCLRfX+IwLiDyK3LegSuXIxPE7R4KH42KRCuERSO5Lc82NNbkS0I8TUfuy6NkezRNR1NL
aULL02uS7A3qALjGpyaYli1PFtkoSt+w9czAmAhfcjx5Ey/p/IeGm2TTFj65FxH2DCEuSCyYxrdw
6sI11+idFFbVduqPbrq/OfC3rdiO2E/amIV9kAE80QAmMyrpE1fBCu2IpkJvpC/9qrV6Uzi+b/mI
lQdXGJ2rmHyKszrVKynkJ7ddd9Jv3iaClS6v5ltzRhPESwk1mSe1kQoAfTcqb3WN3EjR8CTHWsvQ
JkSeuL3Yq/r6Y/w8vrksSklumWMCEIEDVVvJm7gb6/tKWdlH+D4lFXQ9sNIwntojEurF1yWZw66S
D2o/eCGIEoN9u2uo2bqZTjvwmgcYPiw+na5EAlSQNAU6vS2fxIrWZIRQhJCTYjw0gT09+MnOWpD1
/n2D1mY6cSJu2JO1J1JUmTPidbKg3j76jwU+A2MPhE25zlh/rO19p8Xj6JPTANKf1N/OiOkE04ut
Gyen57Xp/A3GKE7JlEEtXTUQmJ1hv2nf4B3dWxjF/fJK9jExfce/g7B/u0RwUoSYGQmkYELS1aNM
VKAEGBtGFQzcuImz91OvUE9yDTjcEZCsco4ORdzlvSng6PsGrjeUAUgvdX3qgj2jRze8gHJ594fT
i6uF58fQXO0yLZ67gWfvToBocuFpfVnjLiTGf/PfswmzIFBI1Skyt8To+58ulXI6uCSYEyFz9bRm
VhjwomuqwzC7KtN4Ja6nkPs9AP+lfC2Uo8K1fHivdCbrK/ONG5zp0TTnzG+XWUce8Vq5LKYK+MCb
YYRfetbCb3X30Vmw3dYJ+5OgMXaZgeE5e1zk47pPRG9RE8A9m4GAeKVeAsxEul8SFlxtS1na6rkG
FIorgt5XLNtgFUbM0KpcNmCt5aDSRIl1uAJSuGoDEu+KgvAl6SRyvoIl1M2WTgmtrcbjeTxdZjQq
Is+p9OiFbTyc4AxpsQ4kgYQYzH/wTNklLeEXH7DSOaKE8xpEQOBm7gQ+6lLiNYgbxW6JPWxlqPM1
zJ06VZ3dkj6X8XTmn6G7X9gZtpR5o2XoCiA9vArpS3ryKTWPHAmcPO0fu9fNpUVIQJpUh+x3mD0C
k3S5GjS6cqy1BJR91kbDedXDLoqtxR7oImK4ev0jxwvBkKSTraO5u0oJxkXi4rEh7kJs7YY6UXhM
i3iL0gzslV+APCH4kPDMpceasuiAGt2LdsD/SXQ9ehuCBn4N9/xyVBdMV/6DZEPt5iGfhaiPw0cy
h8qBPOupnWFjGYpr5SCGz+nsbuhrq7mEdvsGHFJzyJOLrbBErBtzYwl2golsIyyv/i1/r2Vtu6Ch
/IDJHPiqwCoRtn9rZpf4pCo76hoEwpx6gR9mLkVCjSz/iRZ7H8lMsL1dSg1qScCLEiHCSofafBke
YTEWJxF/95HIP8eaAHWWuhLZc+bSh9pG8ZhE2liQ70OMPP6QGEHY3BZ0wzYbiyCFtph8qY9Rxr1Q
GKEx1R2PTZTjl2+F5umCjBY4OqHXyuOr6BuLyOTlxgCBhgxWRPlOJ2C2FOc+4enqvI3QiGx09Nez
txVT7Qiat7JgH4qIdk4gVbtV2ABV8fhvCCVUSrKRcv0oXHRPYoHBIPbDNyNcYsYxHy+6H5wXaJOo
SAGHOH90D0jsr2oNe0JRYPeWgMaiqnWMwZunupm/Q8Wj1cNCe9Tcgj6DSHoT2F2/sB+XRyNwu/k7
+uxvDZtJf8+ghDvJ0pLMLCMoe6Ju8l9KjYH5ofWTeGQVq5B1e53+epEQ2lzGAfMYuSwTh46OpeAg
kkgONdHQeCs8aoQ+ruVrIl8Rpfb0BYgybO04GMXLP0PjIvpsas/S6A7ixN1JahS7YrVi3NOLR5EM
hvTmMZsjUI0uIw6co6e9+I5bYToThiTNbmCFyg2N52iU1ngs2Pg7IFNL1A/E7vyyfK4dHYbHyVyc
vjj0CrpZ3hoXhGrvDZimipW7WC+zDquc25I8/ZKQQhD27WEPtcB7Wy5IFNKbxJDvwEFVOLANxpSM
wE7gezw1KuaK74YoJKYuIxG32CGn7ODpamLAARUi/6QythbfwN7K51er0bvTObaS5cY2f1jI3Rx0
a7hQAQ2/5cn4dOMmB6fY7SxEkgZm8pqbIsqygIWZ0P0B4BhAuVp4LsoiEAhc/5sIV6vN/Js7UHCr
HUyI+vTJxWk0OzulQn2ovZiKKancvF9JbKR808Q3w09AZ9boUm6h1b4GgFPCw7tpA1M9KzmqXNfp
FsAG4XytRIxyvGgv64Q5DyeEAz386QnWPpVDcBUnuRkusczVOb2XgHK7tQ1BvXP/aiVcbhzMr3h2
9iEdLbiwtN0AYhgclOc2DOW4jlmPU9beH6QxOz/nMrx9/XwpRsn1ai9oDz2/iTqZPQHqINEabPuK
dD0Mqt2hM2UyW0X7R6YcRAYm5edkIvRv2keTWkG0tctxWWQYTmyCS684lpHDFsqidgzLXaPjgDHk
ibFwl+kqTFsoOzo0uxnl2Bw1h9YuxZ37Re6rApLto+J62xraKxuY6osiJQo50QBtyORN80f0Sz1s
xkpsNRjunHTn2MpaBDVbwARIHLa7PoiMyf9XYrj066ZCKGWNM88k9wM+cuBkNHuBmY18GNa26yBC
U66mZQjVQUw/7recBIlSzLmdHc/eyAx3s9zzbKh31r8Zgx8d4JcTiC8eKEg+JiWUNPv/iicglQ+2
Dw2vEVagWvmI6VoC0kfa0Vm1j7iIQnCCDsvU+u4H9C61jxtNx9ru+pq/SolJ4L4E5Eqp67N/ZYxH
Lk3ALE7pS5ZovHkf0T7APsXLvnrMrZyozSos0LcedDLSngzitvmb8RkQQh+tvh0B3TS+4+u/aCDM
XAsTKKb7+1CKDigBb3FLrUpkqh2Wj31SGLGAcsAguHYQanui6EVJUS/wfcMPHXJz72DzPHJMe6OV
NY6Lidp15ZJuxgWRfe05llaGbNQ+D7KmCeRDrjS9Ra6jqYX/hg2ekp3IKcxpQFLOx66TM98UiMaL
Q246ToYI9kczcYj+pfjb/IKUL+PQ9zINTVVjYYE0K2yhJUEaI4vyE0I7TehJEzhemEz9ZT40tLV8
BDXCEqq5kHOzRXS6l/9oDtTM6AnsdnlM0pl70E/41CjEHfmKRLfLtbp36bB6JF5QhDA4LSjxC+LN
u4g2MVvZJ6rOUNVmG1GjXUT8jn1u9HGHwXwucAHIgHJ+ZsJiy72UP5MKMvhansn7RC4TXAVFz+SK
gcH6DMIuSRTEI3T1pSOAEXnjF99/VuZbjRr2FPCFZU3BctuWP6qem9iocsXes94UPWWBUkms8MG6
72+hf/jCoWQ9HYqs848b09e56Nad8HJjmk4WTnMpyE6IFqZGA/7w8Gcvf2C48gRosUQ/wf+CBvTK
BY8wUOVMdWDK8FkdWnAdw2zHHGSlzBcihxodw13tlFCcpUKm6EQwV8MK+xXs8tRttjK/T9oc4N09
vePwb164UZyStTtJStzBVuxqh/J3vl/pXZ6AxYaC7pkuwxQW70EAWfPHHFtPD9cFO+9b2WIYksW9
EDcnABSFzX7SJOHvgeKgtvXtV6Wt87doBaSjSy0H0PMIZYSXnY+efAr9YO7OAUynMWM1y6murRyG
AAyZ2Dz9TEwOv2w5uXk2SRiqCVbYlDY4xAJPVnx3KjeAf8izmQJz0oFlLYCVNrTUo5b24N4LX0XJ
rbsEnpHpjgk0zWkixj6pyKZbzbbH0Jl9Og6WlxFKZKvXngjI+gViinkOwgUC7Rh0LrK3SltBfbgd
GSQVGfqIYRPkMvxXkkltYif6/MKiPyMvEVAR0KMWvntWUP0CAXcT1leKlqu6EHd9Hx/p65fZzKG+
E/tSE4aGTIASmYMKqozBSlChEAUiBdEgGKnrFzsgNZ7ZwC184jnMQeydkiczIgslyEICWslCBrFC
9HTCZWZLrCJnH65klc83gtI2OAKTEmPvLt0ajYkPomwn4gGAud/m8xL6PkLhKwo8/a7n7XGgGrdN
xFlaXXuIkv7efc4y5IH955f0ID1lwWlSQlHq+0SjTXuvFLkKaOOMWn8vtf+JR7qjFXzItc2H/a53
UFZhsxBbKx30QCut0/zT2LZ0QwJo0RIskcIuCWIw1miG0jvygzIbBsCQLsYeMH3eP4+AjopK0Krw
9OIgNBVAWlrP9imnabc0WHPEEcK6r2Ek7nrpb++DtKgJqJ0HrBPAz8OO7c0PURpdMfZLrH+iq10i
wpJJhS8ZWVtlBePVXujCAG12vL8QBPOKPDPmzhnSng1xpS5v2cPDjpH48S0ai5k/40NR0wxlca7N
NR6ub7E68y9+8lM/ljcAE+ZODjLQ17t57c2sVGjjKidlVdNUxyh6FBk60OH7eeIBqn7F6b1FkA/C
Yn1wFLBZBr7u8WESSvbK7pR1+bUvPD4hn76PkZ/rkshT3Pq8pNCFPXC7Vz50MkNyfOdRBUvgWOqA
qEto7Qh9gMTJKDvsKfb3JAyoee22JJMyrdimvCG5xA3EqFidrnHvw7dOtrO+wzf4slms/60Gqgaq
5AOrF71ygzHSi0VRU4TJQT6nSHymTq/R8dp0Pkc6XhPJiYnXBiGTCH96saEY9NFbpARFNbEJr/To
TL7aXr3mYxnA2UzDfbpoJxu9ySJV6K9rXoSO7RtBvQ1htvfUmgRIBQgIWwM2qvNYLEgxdk4EQMhW
9RIa/pd/ITzrtAfL1Css/z83+OfsB6vNo4oOc8m/l3+XFOO87jKS0jsHu0XJz+QDu7HZyfHgE+7o
gIbzzNbRsGmUmx36n/fckDm6F1Iwp7qi8xw1ViFc0+ZNmiXcAo7464XMHVvwNfTJtK4JA0jeKgBz
juYrz/i86JtKP0Zs4B0+03ydeHRNZch2y0dLV4wSj0pm/n+CpKvX5jD2pB2a6ZDytVxzgwEFp2Ht
D2WfQeP3MOTqo10tzfu/OxBHrolNUtoIkAh+X3OeGcpAtGl2/t3juGDG5zAv2qdQWEI3TtSmspL+
a79CstDJ7mfxJ3MrC8Wt9j+EJx4AHnMvZQHSPsLHjic3JM22zmAq01x1oSrWY5/nublPkIeVL0p7
ezZRhk/pD8aWQ9U5G7sCbOiBoZ6EI48bdEAdUaEuSZVZkM+d14JgC+9OwXDBNvVnEGXbeARdTgKW
Ado8SYCYRz5fLFxHC8MIHh01Tzz8Aiz1JZs3rpU3d870cvvFzF6AeMV8ZNYrblI0yP5EJvglbaAG
zsuZYWDThfPaf6RZ5BKw1vYY17G88JoMlVCi9WFJ5qAU62NOYo5V9cxRTmjIR5HxsAO+yDZVfB6L
rbyY+X3IpJU4dO68JMDqU6TrvGi+l5FLCv+3Z0Anr0SWh7SUt7o86CJu1pRpVBCnKQ9uaFU4z3Gt
uJGwtBm+44RiinNT2ggyVN7b/RLhrFBkgCQHZ+0RybGV+Y5coUM7JlYDPv4xjhvfOc8pW3DiFP4b
w5Gn+jvf9yhmmegt005td9HLvX/g3JEnCOIPYLidKo0Kh8pN/cyJqxdJvNtEc616s4eNpWZ4tEKU
9uExn2psedrtRx6Ni1BLL1v/3Iy1JQb1RX6HEu2RZCFOQNH86s1lYeirOSn51IpC2OpYa68gXe7Y
Rw3Vzo6xjCvoCNeXiZprj7op0iJxLz+5xi+YB2JGKtZSBq9tOwuuo0ogz3mJwjtZCkxouThQqXX1
uiWDZkaWEWblOCf2hnTACktiTJDmDUUteualEAFUqNgt3EBZFcBBJjOfzD+v2jCO/pDsRtKIqgVC
i1Kuox1JxLdE2OnNeL3Ogm06Q22uNpsu8tpmJA5Pj0QzodktEtNhXPA7QsPufYp32/vabrtAiekA
ckI2w1N0MabD3NZMBRn9UmiECRrnxH/yxT/96lxHfknEr7semoOdHnLd2XqXPr0k7bVWWpuf7pse
krFVTxzKyoOI2ZRvTs+sXfLRS9jFfqoj65a98+fJrKnCjR3BrU/2ZP5EhomDT7pPFtIReM1vylDC
NIaDg2hCtEIZF5ORm8PDeEDsTQKnSagyntRAfpL0PtvZK5MTKLyTczU5zp4RWx5jEApsrDTNVRFm
yYIjhvUQuye/7Xl4aKH1Tk19j2ra9V2cKybP+n2fYQffIdBjB3nYIJdGlFLxAuYl/85LT7e0mI2G
S2oXfpnBEJbl/BPBzvv49U50R4CTQb3E5Ew3hnLHSiNLBCDUCYzMPiDDPzNIkT1LqnsPToCsafWs
xa/+RABExSnDGzZsxsTelr8Dg9sPgdlUafyJ7JuktM+GGjxfRvEv3eEw1EWvfwzLYofo97jFCw+A
ZaugUyvuzVnu4LC4VPL16iIM2sFLHMtEgaCheVDA71NrjayNeeKF2td4e13WPwrGPTympaT5TI0M
Qp2aBvZRpQUN4eNiNVrKZICVLZGs1V4FYyhQ5ylyeAl4ahXqi4iDrKtUNCmhQ4MnNE1/aCylUtJ7
ligyiTSYnYtnyM8PW3Z5k+j70CFkmYL9GBW8QoYf3HmXYUbsaaqyNY7CIsE7LANIbvTLdGIpMREe
+R3EnxCvALcfnESZcYTdAUFujdu9Dkg4r5sqH45sLI4b8b6VqL/yVdS0KRgPn24ku+pA9kpolWfo
5rhs6VuF68beHBdLdyDp13R6GGMrKWTPKyOxsX9g/Rs04PQb1kR8qcDfo5JV1g5ik6751bO1SUZN
fwUgzStJMxiaWK8JsPSvd4SV42JpF5mWHN5iUWFZqmkFwJwn1mr5IMj7BUWqLY9imbcy0RSVhB21
Uzxhm3tMDAcX+dqMVw23hu/xHe6yohyLpsvxRDUvBkN7YRJ0VuUMT6EMfEHnU4lkXJq23GpfFzmN
7iFBKa2/IKEbfCHFc+b+h1ogOCqEeuw8CYYAqU5+Gw7+WVQ737cTjNufztaX6zsbYd3KZr4rp7Q8
MO1ZREdJM79GIHXANbTVlgQVyyKdGvype1/eCnHf6IaCQVyGalJJzZ8usKo8WoUu0vM1Y4DzerRc
C8UEZX/8OXpJgDaQlpOY1TYaVJOLbm6hyLUBUgCCVxkPrYqZQQxE/FDqKmXaj4nHzDHzLPvA4JGy
x2MBX5/EjHin0Av5t/RgaELxon9yC/LT8tVtbo2lb9DOxVpWyjugqs4BbAB6HoceKX24bsJCM3in
vfFbm3i8pF2c4GSKOG/SjGJcVNv++ig0VRcZkQr4Kobtso5pZDp3t/Q6mQmMGGvbbt+SH71M0sBV
yorlKxvWVsAZYj+VV3RG4cOaxi/GrjjfVtShUvfJej5OoPz7qg1YWyc3Hdn094FaeZ9jvy3noqaI
2SVeBwaZacFORsI7aTkLS9iARAiQ1ciqBYZ/f/enG4MklaJGbtZyRV+WauU0yPrxn3zim0Cg6tFJ
GY0jR1LpfcgElBn7odYN0j5KkNitNJdoly86pkASqxWNEqZJn5KB3aqXRRqVIxLyH3wtnh20ivjp
gIQWh3ceRhEOtZOQWaSbj+1z2DZCfezTDUaXD4tjr3DStZlExzCQ5OBNPMKjhe7luuPNOldWx7th
I/036RuQZSACqSNXejCuuAdg9mEoUE7NT3Oy/0ahCj6J8ig6FCUZDW4mEnzxjD8h00Nedq7tlg5F
UvImXk620Andh4znNSV4OUnof540oqcDKyJwhNZtXYaHrCILrUd3rc6a4GXvYVGOiXAwJelCDFaJ
TLImc1Ug5a4sVfOi6ZQbyl5z7CPBUAM52Q5utCp+Nb+Ukx5t4JHGP2LG/37tVGjNDsptXbtuEubU
LhseJINgKIg1Qr3dX/vor+1p5mkKFnAHFo58WCfRnBwchzk9EtfNOJuHLoangv85uFzyEGrPhHKh
ckDfM4dYTsO3KtAPVCxFEkCaqtNw4E0Gp1CG6lVD4S7q7CqkltpMyV6uHDx2GBX2k/7qjDgmkWP7
9Dn3a6TkhJ45uvyZJ+rNN7bBvvq692rB7ztmYxbbDGqB9HQUNgfi3+zxR7Dt7iJib1HPccXY+URP
bzpPMir9g6cSfAT83gI0FUnTczqQo4zjWsXJS7joCGYCTajkGavCTUzSuxlv/bdd+5Ij7wTn7yo6
iOMucmD+yKHzqipLvO7zdJ1yngko/WlIKEezXW4qx84OWd2Mrw4iwBAh2Ye7/gIR69d1Y/ZECzr2
hNo6aSSNs/PjLubSGMRtIEWL6+UpVboynnIadHmlvKWpqn8Xl/rRXK2uSLSVT9vP4cu4bNjAvuFl
vln8Oltbe0Mt58ABVY0xmoDwn6MxNVZwwiwn/vNcA/6nLfv+wkYBMFojEaTaxGATW0p6mtRPtkgN
nrpCDezuIfiCSMorMBHIToP8aoM4X+s0nb802mlUePZeZLMCfkuACeWxyHR1wMGIYKW7+qE2CmaW
9Aug2HF6iMLe+rY/BXpIecrSGoIxchuC5YRZXIBiYTGiuNY9d6xwLBHEibmp4wfrxkgO4oeB5P5M
o8jMbcmnBPNIV/fAj/2idgixlsKn6DYkLPPKLlf2zbuPHMjNq2Wamn89WueGRo2/6l/1bWybx9kn
VkqSBJT0MgRE8e4Aw08b0Hq71smxnHy4k5bypQ5uewj1PvE8hdt70hUO1JmZYd7he1L0wCxiMASV
q785SRYfZlTXGKEJEuyBf/5Q631EDBC57UjiLmB3UHkyEMlGfZvpb7+zy0v0I+CW0m6x9qssyTQ7
t6nfCTUXtOd9t09vjn030yOkbxRVRZw/lBfduL8aPfYokz0WMYWVujTbFDa5v9zY7IZVpkNI6l2l
agg/oII+h3V+Tkoh1lphK+H2xyUBz5pwqyUqldCKw83VuNoShgzCsWwcRyhzPkAi2uw6XvAdsPo/
UpFQGhGbN83fGk4Mada5drtJGAPoqjUQ2TNRP0rHrdFpDcorkCVpW4nxOGvZzWxGbQkc+uZKfjQh
zqw2mraiRC+Ueue/+m/eY6N0kIjQphTSnGBNlQyvy5oo0nj1iv38L5ih42ywLmP33h6CxAXIROaJ
uypWAoETywz6NH2s1d8nv4LnTlt95wK6ZJM5SLthVhbo26KeoVzrpNusiRrwM1e63hJ9W9zmhteZ
UoE56YzaC0xYlCfmKeyP6YdJwk3Hiy4ReBjoLx3cC9tfOBlTuvSGUKHpM7RK620XnnqDvOt57lTJ
WjR3GtLWxBYdo1+nqqymsOJJxCIQ2Nl11iAC1TG7WwClSB6MgUkf8lqsfoGjOLJ2DKC/ySa4po9B
AF/MrPXlIdfQTNVipxGEbP3Lu1u+OOYM4M6Bg1K6hCsaBawfGCqw/Qyb6PWiZ543kxfjZacFKsc0
QspNRi4lbAX7jgcb/1XhP+001xi1zWa1mle+IMEYwV2SyrpMwSQlT/am9ORmhetHlj3N8/cUq9HZ
U7rdQUlIkaxkVzxYv7rgCTWy+c9ejQBWo3zkeUOgMi5vDw+V2HEN96pvqEgjTdpYyr49ExNJ4i1Y
pdKrII6NW++eQhHpqevIGHdcksKXHr+EdbGUezP/hbj5yjpMZWg0f3EaVUgLju2gUesUFLzAExEb
808D9fkODw1Shu0jwu98tI8Ggxy8fG+bo3bwJBPhtqtj7V1jnKQxfRi35No12rtvkxkOZpKNPylp
4bBndJ47Ng31kXMv5U2leDeAhQspB3CU4GoTMn/l6/zWN3aeNJLppVjkgkBeTojWqbYBwwFq+N0a
y4vC/QGSHQFRDM2KfudAA9G6bjSLhsW2EkVgaaKcpUB73FzWuh+AUATmlHyzHKDIxpzPFE00eX7Y
eNSCad5kvwVo0MUDo95IpTY6I12JEAIQOQdoY6q4nkrcj/u4GjQ/f0FGznKoW1Oric79n9xeRhMF
7wojJxLpO0apXx1QJMGUZRJDvTO9rzz3mj2NDHaKunFEvNTOIiOBIuGZl3gDJKFGQZj6/cKk8Rgo
xbpDOp87O44g127FepGX092HTPpGqoMEsPszCLdK3a4R6w5ITkldnq4DpVGuHYIlXHYFy4G0UrOz
MHnxVukBcus8+fsKzoEf0Csi3oz50+vL5TVhgXev9Ilggf6OYqp/RcN9sgbir3yJ9/HrMp5jXMTR
Vc3jWArOY4N8QJQ5PMzRkctrm6OjicBUCJW5jQJtVxuG0zJy12IsXGxOp7p6xOsvqzS69AM280rs
JX1Y5qZabYETSlp2t2O4Wn50NdsYUHHW7THHNO1OceGUAIGC9MxdedD2lQDkWIUtBLUenqBZGEuG
2N3L5a3YP1qagRVs3VpYBQ0TZD23aPo5tB0D7+O/LLqFDmW9vzETHVM/ZQZah6XPrJVvC6E0Sg/L
dP61O7bnGfbJsRQjHecdivL+xR6TmH70bInGah7GRd1wNlFKPUEKNb/hIYZvvTHvAi1gQzEFS2vH
NXAVMgMd1CJGzI55IwBurTZpv/pBOZsHIImVtKdYg+FoLq0H32PmYuiB14heIvsGZGXBDYndOPCm
3G0t1e6dDABFpl91kr+KkPljKuHB97FqwKQrQRCS/2oQLFTxOcWoQ32eNjtNNDLNfamAv98zXMYl
VtGZn2CEh/ZBLehjvS5EjJQ7y0XSYvJBdx1qtLPmTXoHbjEpKkL4uAR1ZiOsQdGOjosaP/p40biA
LMg7UroAHot/Xu/ygq1tY+OPRGRtwyOm1pxsysbbNlOHLtrEEFkyvyU5Tmay8TaMWZs/LLlzFw9v
wpWIWhSIuFTs6bsfCQ/ZS7gyALh3D9Gdi24LHEyQZ3YH4Cy+IX6B1ygEOo25d8mMmBhl8iQgTXCh
AsScooD8DdOHWPpnRMoYsfBQwFzVuEZkkTkoV8OmQ9iTPWWUWDgFX+kSQB/cTgXV4QPtFQvTOtVc
miXML+we6mhSrn8f2OrB8Vmcefj4Y0bzULZLZrQaVIKvJdOOsqkTEXQhYMFn+aUfNIEZnbviFG0i
H6/aWV0BCudJJkcFS15ZNjrL/hl8pk8m5ASMbr5lizk9Na79oPhDQnZ8+XpDqbABaO0fGgr0WIDG
NnJzs2EUsZE06KD4E7dJbJodfWw917UisI0Lho4akDXAbiYCIFLSwmFtP+TW3Cnq6x4oCtvYe6zo
78mCnzxECEsUXlrDTs/gKgwoYSSRDP19ee17gg0vUB3DN8HM3CBNEuhHcq+fLaC8kK4nwonWwbuw
89MMjNvKyERPTDXw0pNarvUicP3D7UVCJvqhTV9hmHn0jeCS5sRnEoOH9vOD1FXGj446+oGg/nRD
ntpFraN1ZN40Zq2OyLT2nF2Zro+UTyfQ0HNMcWg/WA295aGC5mlzfBLrGor4uWqxYK5asDVZa5NO
cPucnf7LdPSM0aqF/FNi86Yiv19SBY6AQ+5nKvkTavhHOUvhb6IhzTZRHZU7H51OsU0gs4OHNOGW
BGt1jNQkXGwj2tl+rFsW/Mxgagd9ycecMcMzFVtn6wrpL5nCXXCbcRJaOBgJlqC7Fjj6LB4v7DOp
oy8LcaXrTtwMv4V+Ko1efeiiNdCd2ijF6plXpKvT3n/gHLbsdXJ1BvfAKNrMpkrjtWXNQsxnG1lD
zi5opMg+eHp03gKp0uPO9Svs2zOnk0nnGuyy2dXJasWKdN9C81CMqDQ7kRqNTVatMYjLl02l16uG
TgnFh5sZXpWkDDR7uChncvHm7gkAjbhTjMKl9QrqieAMHM1YLq9SEo7LL+UuvTNpIKE31cCUSFss
QsxdxXNKsKGXVYRS4mRLuyKlOuE1aFXCEgAAd/0QR5f71qmc/bKr/XsQ4EQ0pXn1MldYt7qBhYsp
X/XwLOt00gjb0Y2ZJH6gavFLa1lzw4MHB+yXhQwgaCGqH/XEs8nWoH6RvIKKyMriLYuioNEHD1Ao
KSn2fluFI7lqOZlNj8s4hQ5EQJ+m+z8B+/3uzoD+10YCl87dTiQ3EIPzqUqWfUIEQw6au1XWY8b4
naYaK+E3k5Ne1Ocs5D+f9FbCL2iGfS0g9fCyl4zpC+xh4YE53/UgIhhmWHw5yZl6UMHbRMcU/bR0
oENu5M651n6ngX2BVL5NW5wO5LBtzvvmFLaU73XnB8cifH+lW4DHbnCCsY1dD+pM6h6UDiRtem8P
GuEgjdYcY8YQFYuz9SO5w1L+a/DOsOwB+uQqtEGDMT3Zh0BDhqO16YP+exVpGFqwx2QmCgoHdbRg
91v/zLLycBgli/hGBA8mXlS1XeiJRdZXBp3tT/DaCdgZXGFw19Ery5paPZq8rKiJpW0ao02MgKsW
QjIAMMLGJzPpdBL5xrkDRnBLQxkuF7xMy0kj8/J042n8bTMPHcbGdPbBSkoFybV3NGh5/+Y4QhBR
YVzjgBUrCYOp8PU4EYqzMxE7Nnty5MsPwIaQL4BrNrPLELeqDNwdmjHgUk5rwK+A2SKi/F879Ghk
le6jGDcjJ+Fpt2qTD7TUmvL09xlet9u12g5gmUw9miR+c/WRa//YDkq7oJ1lLeOfT/PMQ/C42F8y
gO25mXd01PU68ituKsw3Vqo2Y1kJ+xOTfcEms3RLggCn6qWOKcQltO+JRhWbP+H94/jsQQJn7tox
3n0nc0m7505sFaVq/17QR9Ua/6TgdWswHfzyYqp/rWBTB3MsfoyL1v++HptUXRK2HngHZSKWEaqN
MfDch+jOp+OceVUyuwitTrsDZLrADcee3FWB1a9qbLq4adAfrGmXAvx3kvoX8jnucvqqGo/u74Fi
z/uHGAqsUbYjlwmqsKZsYnXunAyMsLNgUZapufaTieF3XbLTuTgaIormFFnU27dHu9t7IWqPKdc/
j4kUkWpe/nWRnZBDonw8DZohTppPaWOKq4GfFc0FG5E45HhITM5h71e+wPhWgz0sIBKrwMPOuy40
Wa9cVcXZ85bFc5mPcptTX9QIGfoIUNPuntKSLdEcaI0w/fVlkjogKi8qPgFnovnM+0322mwiwzhp
qcXrJ0g7JJLpGIrB5JL2JVxtBJoADWgA7SF28Wu84uZqM3+GfFeUK9kNh38Jzs5DUHBW64dmjrLF
Cz1blJtloUI8Ew53QwBbT73XMX9HjqDWnN5rWxnKT/SXFW9VDNDM+FNbRWyWMTP29jiO/Njtct26
fThZNkItj8COkEgl/Qmr69c2kKSoMT8/DtVEZqD5DVptu52fby8bFDZC5nLol05Yf6H75GoomgRZ
nEA9IW7DFOuqESBah13Q+nlPRBxjp0HXwxiefSKuM7NRF9mCKWIaeZkdk4tm1lTTl3UnSrYeaHXc
WOI//dfVuAEjZsGKPQK6P5eXhCq3q3RSx5kTOZ2emGBFUw5VjfkPR2l3lphvl96VFClvNDWjq2+N
u5y3o4ECLbLqO0D8C/eu36OS+MNCZS6h0L2HTYiMgf7JCDYlTuNjRJdNvuS+ukvJQErdS+No8tSL
XdVRvVxUMs2HUHdnffbB0q4QZO2wmFhVC1prxz8+04bdMH5CquGqAIC9r9Cu0/psacqsAzPfzOVa
SdQ/OxMrZc32p+YUQWzhZQm5Znp+aRgIUbV/tEBvjSTIMlzXUFklbrG4e9KGcqpMNSSKRqfHCuy8
2/UwKQmJgyNw73Hocs71byQLCrw/+3mJDa0VNDDNUqH7y8Z67SknQj0B9Z14mXC0bz1rUI7f/1Jq
40ocRc5WAzte1zQ9GvehPJ1ORUzZA8SdEty8GfCQwAsECjaOKt3sfJU/qawPvbvTTvkqKPnd2ROz
W9d5U5bkJW1kkACEhs2pIkA6baH9pbXuz1Zjte0PaKAUTHBRufmg2IY5iHbSKqGDGK7Bej6pICrm
ylE9OccIPddh+gEvM8lCNrSXpd6VygHQaLdnF7oQciX9GenS9A1B2UXmkWGaSwZsPRH3+rjNxa9Q
fRMu/8/b83NsfIhpoJdFgJUMjIZkzSJaIm77RZNNJggo4YOyDqCzQvpAdQ2nLpXVwxd4U1bDFk4o
yUlk+B363y59douIyGPNuwA7pFAuxMpbibgPqmrxGnLUA1fuXUgALpuhAdZxDbtzbYU7NJ1gdm7C
+x6qQievPFjDeiop2LT2byjhv0kQ9TwJqukYMQeN1AFBA5Ij8u1xgGoB4gYFJ22ENQH+ylSLEzBq
CXb/kz/wzqkiZsYzkWgXs3oK2njQuoB2dAagxeemQ4Ie9/jdcxzVxZdLeuTp6ytUFXBsKvWGmRyW
MpCkyGLpsYlWE8aU4E7gfrEB4IrgTDeZcUC9TwLwtHdkOkF9ZlYFFfGx+P0ZSlzcJOyF8GD4/rSL
ynPcvWLU0fDm7DCeKdAIeKGv/qSq6cyXqERlmSiDLhlLub8oox7TaZDmtOAdvYDaAT1m35SSjfcN
DCCcNEozKcrRRMzw+apl/5HkhUNw0dKfJ/9CgLJnSiyp6bvXklOTp5jWSIzxD+hHp07TdfCF77C3
J7FQvlDNqZK2yfyowjK9b3rl2VSYNFhaAGPrcbUyWXdf3p0ay4GmyFXpzRRIZ5pHnBJOEZmADiap
i391QK4W7gVcrtdRfqdeVJiqlf1NXCAm5KZlKBeEf0JLuFxuM1MCxQMGJ0m3qmrzaSt+SjO5N2SO
kYvhnoKzSIqB3+J3tjGJvBfbMMjI5pBXopFTBD/f1Ml3IdGpCT0VXfPJjHHlp0nQ/NcppZ6HOwlC
u8OyuAOF4I0E/8NM5w3ZJwo0N+ie8mL6sojDEvvOK0WujkIEXcVvHsgZFkILmofs0AZkEGqT+Dpo
Zk/zLLbEW4Qh/T1sd386xS4U6oe+HErMtBCHpQpT9/lZm9ORdlfmM17Zt3fkuXB/y+QC1f7vhFLu
U1yndX8NEniFXHmQZ13yiIsyp+1o1QdHdtypGruXJvDjziMYziZR1SKgkNafLtRNmyKWwUBVQT1N
IZq5cFw69BxmIy44JBNBFL0q3qngIdJ9VnfiwW6jHIkvLpYa8nAiXPy7dqlTtqehjv9t4kRT3x+g
9o6FRJVTZhai37sMvfm/RdtWVBdIw3iYHHIr9eCHRl/R45BcNYVJYiYZl3EtI7l2nPIpTuOnL+Zq
UTJy8JaQC0VCKUqkC3bErQG30v3zBEzPzJTgNgOo3Jf9JVlzmyRTpE+JJ1XNu7o2Elw5rXK8QZq8
zTQ9jFQOOWIqGw605ibT7YUbj7xH7LufKxRUQqrRY49ea/A8rX2Xy2aTt9qKiQEqaPoRmV43QJjB
Qy2QqBJiP2SVzlOumvnwXvJbKeAp2DWNh+9J2Dfkx9P+oQHJeTUDaZvwUrthHakC6R/EVQW5ceD9
0uaXxSThxpiu0Yu4D3bAmncVXvSoOC0lo1ayT6ifsb8u/xHbs8T78oblob/i6Yyk4fgT3it5XKvJ
1BAt0pUlQr4T1ZXTG128OpcoCrJoe+4hNeZrz8wTQBNo8syZFgZSmHjpsGv+C3tt6lxXHTIv4Qop
JthbmarZkck4lqA8n5nbtkw1h/L8JDVu6PoQgR6DmcqSQpo8lnL6/vZEbTmGpwMbFBnvSpcsZ18B
RD3uLA1JpME4qPu7xbVSqnoagWeH/28tB0U2Qj7CNrTbPA2x4EUYBN+DoNJd8MA551EKMu34h0uU
3+AOwElY7XdDqQ7H1mOx2XW/m79ybwIC9h6p0/5TCUFziMITnlLpWVWKpH8GpFBIptPd1DO60SCX
U8ojnb/mPM1HQHjfF3rSzGRBviyqxQ6ijyoUJuEie70mujHWyw2WmxwGNxZH+xoQWm9DT1G7anSl
NqN4TYR/gOdOhDm8j6Dps2dLKVguxpFz2MI7ujBqF4WzLWMBd8QTe0AgBs9w6s9McIWFLd1Sj+wG
VfwwF92WwF74sOWtJDcQnqlEVVe3l7FwW2LJhZKEX3w5rDEVz4XcXPkZpmhvVK4xJtleldImFXa2
EczG/ogFtzclir8UlvIJt1knvOGOKJ80vk2lg/7rd0svdb5t4W5AYTB+RY0Z2G+JB8fBxRWAasDF
/JjkwlO9HHNap5I2+2Zlnrxit6ZXNvBGyb0jkjOzPlAKIJOFMEWDBtRQfg2uSOJquTrqAprtuPd4
4yAoBaPUNm1OHQppZcJ1dYeWG94g1H+wo5TLwHq6tmbB6WWKldYuBFrObe82G4QMHqppEslLi2KC
em0+UqaD0cC42H3H6tMmXzIKkY84Nje1gQuYd3VsnS4SZrktr7R8GIit2oidTdspkqGLiu2safrW
aYootQfvyK9hSQSFzP1L1J9K6F4Y58b2b770GddD0ZFb2atI7G5pUZLmeGsoOY14i5njQETjxnjO
IKFtDpB3fHzNrXmiPsFpqde1sbYNvov2laZ68JLoS+u3cQ17PyF7Yzl4hF9Ctou8vZH5JTkshixb
PR79H4Ms6gFEDyODGeuwLRGHCLiIyY1g1/eCdprsHysMk1/rh3VGfa3IOJpyS6nBSJJ/572KI6aP
rg7Ub1OHCuFXQr2VtmyHRYdN570yqCH28p2he4OZU7mIgDmo/GWnG16xx6HlrgPSjugE0PBX65eW
1IiHnRppGCcrfYBoAURL+eyPUzmMTQblQg0tkK+U2lFtmCvtCh3kQRM9f/szwq+FWIKmo5bGtkX6
RG5U6pUtc2GVZk/xlF4OAHyrUgLJ7N0BI3dtr3JHdaOz/Q/oeEwSfjjrIZ3Jany1wBJTOMThKibR
CuEWmn59y72S8QyrDM3B4F/O/rWWpiA4dOyO/KGvCCq+SwtEl+NlzwE8DxevcZupF0gvSj9RyzIX
ECBqg3EjlJHifZBU+N+QB+23yx0gWhIEB+ZEjakk2IfJaXZETeo4+qygd4DAaOpy376a5J/Hm5Vf
grqjH8tYirOwX/iO1CMf9cTQ1mNa4lA579YAf9Yz7e5Kvak8KQ7fGkz3kx+6Bs6bDkI7f6QSzpwl
BzQbTJtQTZM/tIfDzxcIlIHxDNeAtN/ZYUHiC/gaYRlYb81TfFqHCrVZmooQi3EVo8a7Ye9tX7tI
DAQ1bKEF22lSggEzZCV2cJqJ1JxZFCRdTySlCIJFdGz7qsQpUbuk3imWUDI9GMqZqO97beWO2j5e
//TGwQU8ZUEUeEILi2T8fjgo/TUeCy/5D2MqP10UQ63tWZeIn02vl7BbMB/IUFGeTPTbXDiUwWC5
7kxkdUx2RRWi+NTd8RtWw/htuCKbSV1ztCkM9Jeb95BR0LYFUMoLBbTaU16ZeGxv1Z9cDJMED1km
ws5uYuBoZO1XPKsCkWZ12wh//AK8a1BebHB7Jdun9h3oC2A48CAwSmIsGciPqLacY6q1jpvkhQHT
C/kuoRpzTJEmMX/PjFnfeIL42RzgXHGdExYhbwziDFRgcPhgJ8XGxQ8bU5OhfjFIN8PAiEDpRGV1
IToI0m/STjfXGReTlaM6QnOSZkzi0W9SgIXnjTbH6sAQNAeSd4WAwhh8cCh/gDSqw1D4MXs6ZtEb
e+jrk7XAe4/+M8JWJjeyjUnnmp+uE1fEUoBS+u8eva7PCmhjnBcoWTnBP7W8I0EzBVYayeV00jmH
b3sF7eJczfsUJMescitleT5D8+ccqlHr1Gyo1phiEoJptihHUT/jGqTZ78ULyRWu8PY80vcflziK
8sLkSkQabCIFmYks0mEihBbY0mwL9w6KXd814n1i/p711EXoQcfeARNLiFHKwBefUcxucQaqOMT4
Ror/989hcATFK7KNQaciL+9/y2LOSPxSKlCxL4qdnJx5KeQ1iuf+HxhgdIkxsEp/RPWVaRMct/Oq
9cMqQU+8AC5mVWGSpxoTaWBnPaZofd5OFiDG8u8AkumvFoXfbtlA/VgbIf62cdhYiVXLOs7NJmUL
Cpg1mCMC6ow4QUB+bCmn/ibY8iJ6x/JGD6AeXyCE6J3JwkpcQ3TJZBOPTHeHQa0q+4co8aX3OQPI
eLu9Y23v9g4uFubZOlfgiVzCO1RnhjlmBO2uG65hj2iqrYs6MD7Tm7Q7wLPs7qr3cTZvy5SaJDxr
Ej78pH9Qz/+Ps0x4GmfXmS4KJGZDhTKnvJvEcOz6oy4jHnwTZcEPEcowtgG1LSSVegctvCIOyDOD
EiODEqMlYQ7Kvz+lHJ8PAlzxIkhfuGDSt6Oz3IddrFZlBwI0+r1NCYj94g9lH+7aWZ08NJuNxocH
gP4+UZBDbmXcwfmBCLMbWAZRUYDtoPWwjDPLpG5mbxNcWlBT2k/4eFU1D4P6RQ0aJqCOjQKiYzmw
HZtEUzNjoZpNURTz8yTZ1O75LqsSMnclDqyqYPJqRHQYU6OsQEdzhxb7w04fcqQLXCL1s1YiVmnh
wzSMg+vwqL/D6JBGBvBq6/uBU8qEqZ5/144IkYRp/6+894MxOIT0Wlbbe+QYVf9hs5OEZFXb1euc
oXEdXYbbmR/a+deQQ4I1KXeZXnjBNesyviz7GrMdj7CjKjFE8t5coCpj9IfFM4dpp8sAIxfZUHER
0EpXEL+KfrjtT1KQpiA4OKupMQEnjH3kKR3YXxGE58OUxOGnoYe9wQWl54YTDcf8Yjkb0pCjBfaT
lIYwqprbc3j2pL6DhJiq5rBbGu8WrRtd0tnlJGhbyQ8S/4Pb5eSs2xemi7i5Ruv84N3qFo0aiWsn
CDX270cDSNVjxJ16PAA/17G7swZBTbLz+ntZFW9+DSS/RtqKTkxZdOc8wQDbKKoadJO6gyBGqrpO
X3QPwAK8ZZ51Awc6H72trnAbJPGHcQAAtLvabtIDrPWknrBPLWZ02tIsBbXcRVvqhuaoy9oo4SFk
c2ElUVzqk+ChHmgUEoZzZ9LptqXxd/Auq0Tpu/jft+F8JnD+QteDDTyKrvVWLPK99UTX5//QDJTD
F4xKmiRcp2EGa2Tad8tXG/AkOHUryfOzlr1X7cTADUKiBvL8nOjbz4DHUa5+3TUqhQ3PtZrILkeL
fYl3T8g0X6J+bFpolPv094ZmmLtFTpv0yuY37b5/gOKPXAqtdW2SMalkg/XaSW0X0DD/YLcPjrLH
8aXXHr//F52cxxO1dBL20FXm8qdMoh1BYp31HPNgpyZorEiv+s9fHtoyBHrksUrMCHHggIyu0qpU
DX/wmLpQahsgMmVwoU+JgTkDtsO+CQPv4U3edil36InqStU2n6BZ/DgL/0ipHRy4tVFt3bJBqukL
KuMXGv2MwrRtS5mQKy0CRI8fOdAP7Rk+8SbRLrc8AJsRoUPosn9kGu9gT9XcjC77MdQKEjMbFbDH
3yJn3tafI1y+V4lxGv5CQVX4UDnlR7pCEIel5na9dVGmQah+iNJ4Lu/buFJ0sr7Q7pWo0s3TUCG0
1QKbzx+58iEdMdLa5XbPoa9xWjz47Kf7W5nNK1sLXYiHyetinsAF9MAfM2xnh5nHrKR+HUkpXCj6
Du4jSv+yoe4+aES9v3czjPJi4gGuvEF2WgGKo5bQLHPKsMek+B06ZpUjdX8YtKS2Wr34nu7UonVi
7wCdjas7lkOpgfz7lteNs/lrrHMeBAVAfBc4WQr8ULYQ02kZ/fCIp7GPgWr40ev1F9Ddqj66kpvH
YBxd3koM2uQWYDPA9MAmNnVqxyc+Uo/bjr46MnGD/qYUwytpiBcfOcZdlIydAuOXyLiDfy/ljQJX
SuR3jU8o9AsPkDcazy52SikO1rONE8PDkrJ+0c9VnxIG15p88LCg24Wr3WygAP0RFXtQiE2opHpX
TjtmZn2Re8Sw5YmwaK9RZf8H7aTLlkcw3QKk82E2vRjIKew6tmhHNx13W6grqoZgcHyU872x7725
fDEsM5UGdIaTtGQzpz8puXaolUp6dZfldaY2DuUUh7/nbDMN7GXllwlBQbaXnO80d0Ab0zG+xj1C
5kIinJ8SeJbu3Fd97yCcww89mqZcn6qAZXH79Tam7fahbceR/J/lJY860xv+mTfvt7PhIQJLigwY
3MY4cGEbYaJfQ0OEjrDo+UiavIHA6bjEI8kum8YXSPNdZt7NsesLPnLE0DySEkBnCvgkmPso7EOl
oW3m4HCR0s/+N0hmBybKsqG3qVo6qs/0yGeA6t0bCYZ05M5Oi1Ff6vH54N6diLdup0NmhbpcFZTZ
yD0h5HZ6AvDWmYURt91+KeJHkZZxPBwJEYay7lbr6CFcbI4YcI5vCTGmHkUggd6fVvlak02+Mz9r
LQtN+RNIr84abSN0XuXZdcbuZFC2r90ZQqj4pWIiC0mV1zGbVytWGQW4HvOSUfEGNvx9tycmy6RT
sHkHzamDP7V+NyQBF79NCDthnncKjsVzNruFt+AT/E3RrbL2DhTylT4iYWzA4VmM/WeosoDNgEfj
KZU6vYC0srUdunXaUsUS2/bYxLjVm9xKRh8mOg3qTS/IXE0iFS0/RUMViSSIdo7I+ixJN+gASNHb
CWCglo81owQ6eQ371o/k7UzWlGzwlLOV+4t30zDOHfMFXKrigBlYMuCrfCxvq2lW5D77gJqtan6+
XPwOhJ/3CxGiH9Re1DVHzIldRSvk9JU7D+I/RyNrbOFHtrd2F/h6pP9Mh5DOzE2+DLQZ716D14OB
Gdue0Kt0c5+hFDndRlvWVAvR6P7G3qFtwqu+SeDlV6rGFytgbxBZhh/OnfO+d4RNiUUztPNWBAX1
qzTVScx4g0AOmJYkrjCRZpJxG0cUul1gZJX2BQVhfPTchkKX+UsEJ+g5fxuMl7a0IyIkPESQeCwb
gUfk1Lu3bBeeHuqo+yD4xYFazHMFn1dVEPreX8uioO0zdTH1eP7NNn2aLpkEKy4jLzZmCq+woCAj
q9Etr38YckUg6HVPazfmvswCM8O+RBNijXnz3Vw1X1h1fuxI+wHe0v6vZGMnGTN6H/nn5JdYnbrV
rDSghh2b+RNHcZjcEx4IB2zyb1gvnfzl5/ZrHwmmF42ie8bxkZP+CbkiEeu5+E1i1bDfc6Uj/Ofk
5+C3anKYGkRM3nx0GGmL7OABlqLzzB2zCIS3ENovWF/GR4+a+CTqk/enog1iSidwX5+qVmyK9qK3
GzsyLPgZn78wr+vNQffJL9daG9yGbiL/IeYj/DaVnKhsTgj41wougcv32/k4g/QtlYzaq68EDgb4
UW/wi0SSVtmS7a0CmNvfvl7VeumAVRmMkFgKkL5HfRoj7Dy6fGW7XI5XrY+p3kA7KO5SdyHEURca
P6Dq2EvzSAi8dgFnfxah0M8nAFs+nJpyq+ODi2YtJY/J6BEKyddyeD3l4gPB6s12Z6ggSJg84SwU
9m4SHgmfMN6mNGa8o/3bHZxScvTG5nRtez0xbBV0muFNwvrrUvTPP7rpRCi+0LdfyVnsd3ku1jR/
YhyVCAZz1Sv6mlH+w2TfIw+Nwno0vKBe9PNXXenbupwyFe89g+XK6uJaHFKvmCB3XMTpxmyNFBsg
SvlzRMzPuiMxg2f1ZATKRrX1Hc7lh+gy4uH588sCRZBycSskIzEuOjjxSlVNcNvrvovhG2JafDis
7H/QcHG87v8BXF1+c9GsLUPeBcjM/YkmB02dDn9EKCx8vvBUe35Bw2jtuRZ4gnsXBQAMbBKKVWiX
JQIqJqv0t/lagSbpUf2oXRQw+z2rLzEPLU4NhGua/SZ91m6CLhMAGq+vRQTuGkmCjxJF9t1uuQjw
G5hiuoYhGi8SdOxOQm8XC7X0Gjk3omvzq94SvZnXfKppnON5sv7ClBNwRHfYh3hl4/3ipeGGen+3
qNLr8qBhmFtDpzdfqYqES4TGPLbBROFlktx5iZl6HFoIx6hJFlRpezLbFe4nJIKfOzcOPi06TWbD
7vboQ7zLI7WeY8S3g7YHdn56DcJfvtq5UqUfTNvSNyGBpwXSXlWv4N7oIkjMLPUSLTtPpoDFeX1T
1tJsXwO6MGFEYjcHZIb2v63cQgaWbUQbwCTxeVu0aYLUlSB/958MOKt8iHbPEh3s6quZnTV5EmCu
rndd2Ct45wLoVW+gysI6PZ3ZphivpLjDnZ4CSFdmNwzcHrl0fD/7pftFliHzYXXARNRIiFAxXe4V
AnPtaKarFiMa2upjDmKREVz1urBwNwxA301G75Bpg/N3M51psIh3dfPAL9+N3a2THjBQ8suSmlMX
Xnpea/Y6eSizSnm++bZqSZistt9lxblp0vyW+IP3v3V81yOcWhwmcGcU89w5WrxdBG7vzLaLpkwi
uzSRm1knyan7TeIdZssIBoi2JucVJazcRq8ZnyThEGptjc06eCJ0JOqxVdZiByumN2oyTBpjmQ/c
lDMuDjQvCkER3Sin29rjkfRRqxQV0xiZmd03Aszf1Js/cWpliwVDXQfVMhfzTaoEnNZai5MPi3bC
cb6FAP2eoWDHcObDjBGdBf7kx7j7xMG0SEcjkUpb77MUNLYFqAKv145RUgr+zgyAMfYjqSW4Ss+u
LhIlTHtZ4Wi1B5RbttB/TBTjjWuCiuJat4YGHKtJrLcMVdhdUx57weDNkl3l61VVeyDteZ4WJR0F
esnEjjBazw5EnXuB6x6M92YAYsxSscdC9IAvOzEgfmMErccxKzJLxeAZFnEVZDRFzqnNaqJ3eGQm
pAfapmXAEsCplEvwgccXQ5Oi4Z3P8RkODDRIyULLbXHVy1ccNXpyauxkcL3Vd6aP/nJUhlzkUFeQ
JK1zEqKv50E9UmabaYzImPXoLiN2q5sOFwiF1FlL96WQWN2rKkYiXnguAg/qTYRM7QGb0eVCF+zi
xL4OcWQr/WiVTxmA/24V2GeakKmRqrTv16vUNuvrpxIiKel/OXpkUOVpe3hnMT2lSp+WKiYyApE9
ScCmYcsYeRNETHdVHh7mcWWfucPN6AI3A6dW8Aoy0Vo75UVcPG6EjSnXlKPQ1nbZ6zhjPT35iquG
hgQmcS1/psUNBXeBLAM2lzGBDODSni79cKiikMnvBAuJDgnpkcq5TJBh2tUjhoIf0StPLGUxpalX
YFFDEx3Sog6kgY0Y1N6d6sqy0Fw+1nu1iu1G7yVFX+kp42QNzKpMOjIpoQcKuLsy7SkdkDifZB94
XOB7W7Ar1+oBaXK+i/kjwa5Fzj75LRTpkJ979gA3uORtLoEflqBTU+BfP0ADPHY6GnVN/1ZKjLRl
3+fdsPfjJqusBbBvsoeBmB4TUPSmxMk+pX/nNn4Gt420UsFZvGSCXpmMhFUCR86OkQRi6TJTw8XN
d7A6xYrIYzcZMsicQ3J4LDKFFndMB3t5+dpELcK2H0leuKZXtCJYDtXmHi+AnboiteQ5o+O22QY4
dHXdqmHjfnVSwcY+YEr5FQlwqzrUSJ5EFhLp+EcZRI7e3kytY2Qao56jH18jvvDQ2KAceIgmuBVc
nFLN5tCCG3/jn/xdqHOySI6gnJc5sWsmPe72bOHV1BP1vU9PUdVeKiAgr1qK+xXudHdl04TxJQMi
qnZKrzYvRWJ3vTP92jEYK6Gxej4vW+QJp0pR5lYdxajIJsk+WbqWcVYQX8l8EvT8co6eT54qNGpl
qsI6NSw9hO4gND9Web/jKYQ1RTbZLyiVQIA+LP9AmAE+wZY9rJEPuM/UjzRnMq/OtqWwT4QJdcbA
3DV/BaxH0KCODyu93Yy7TQT9olwOGNgUZXZjZio4IsiU7YmwlBbbT1OoECDreGAjO/bKqt1T/A9I
VMcrIYGGRu6qM9Nsm6Vq2i7p1QijFfMrQLtENB3LheXGui08PQ9FjbzRRCvwNzgWZw0rWh0bjWHk
6CjwDr+aRzaxKWNnu1ezhK8MBdXhwA9bKmaZ246j5E3+U2e28uMU3ntxRQuWG2UYuvAK3rMalkL0
/8PN2aqnvQpI0ZrdF0Ik+99wKgC1cQ89wlaQkWeLseDSTgNpSJErCEVQrPCju5Mbr06ucHMM+GDv
LLXVYYKiCTBlCGZGdDvBaZCoYWhkryFmCX2Dr3lara6bt8ZI+RlKyZeyz8gVdebZXLbZf/Hi1ECk
tlSFi09Msl3qQzXV3nO+uE7FeoBe7gdutjDWfS+HAFY3hRB5vaTXwD1qtxckTP6hsxorpBY5yDhd
ve+v1TAC3K/nNhJ7sG+wC47C9zFoV+l93RVGBiWpc0njuuBxy1FzjkUqR1plo9sMDPH7zBvQbCu/
xfg3tk48+jYRMsqlf9FafJI+Hl2XnsDRuv60OkYlHNmbHJ7gDQsHiREzKI51st1XrlrWYIWpg5a6
qcOA8l+ip62DVYhWRdvN6/87hJ2eFQw8DHM3atSrFs/Q1tLNhHVopzr+Bg7B8obE2Df5uXtMuVFk
dB8Zjj1p1Z2c205ZJF5hnOHa0eqJC4RGUF5ZzQI8tCvDW2a3YLctesMJnlJWq5DnWP2hTb4vjH47
luJR1mTZL0yo/vO+D1izGW74nd+vKh/mojeoypBtAkEg21U0soEbsHbIgFx7of5p8C7txZNvYpxR
EWPuF8oQh8USOTDRt7Z1Sdf4R8SyjSYzswiIxZKqzjULaJF4jyQOMc2srfzWXYyF81iqMjZ9yG64
mVAXJ/NoWfmLkdlccCpeNr2wz0u1i9NbQ7hXApAdrUInKMy6rZgQC5a+5Zcy/k/G4w0vDW5l1E6I
fiuseCKfSoGItUQI9wOJa5k3qHdYBf3ynCtKrTYSUx9Hvt+jzNPQ9r8jC94o7YstH0mFNgT60Zja
tSo+IkRLXVO+EdJP8h70eLVXmbb4GaYJH8y2ktA8x3KoXqpNyQboh0wiLsoOnWAA/WKR3V+6t9K1
PCAVRzCYzU0i4phwbEmTHbN5kz3SL4nSnHt7JhK9SeFrkoKwkr+IlTDYvzmYNMNoeIICiY64Bex8
O+zCZiFxuHtwiNOEvyBJe6HfMC8Vlyvtmii2twXcBbFW6kBgFa1SWQXWRn1PBuWfiZPDYKr6opfR
9+LhKWGt4QmrO2jcah28A2JJw7nPjlFY4O8MC8wlHhuFZ6lxhsdYC3tzdRURJmOyJ+MLBhrTj+tR
sUFlzcb1yPVs4nHxWyaGpBIjQM0zLKWgvA19Mp6rhkMBHHDIQV0lxkHbd4n35gSehfx/RpGW8HUZ
oUk2srybT6X55UcaXXBBsYqxtrSwDqlhkto0mfUJCF8L3OaNpTJS7tqOvid4Em1AwuD0DU5vST3G
qqQ731A3WV7zwC4gu/Xxxdja1mjrh0EnxYEe2T4O9xH5v/qi3fhTUzvk4n7lPOOen6AGPjsgUyQF
Jt4Yr5/yTVh4UmMGUGv1GmAZb0erAgk/Da9hyahe133aO73BYMlgBAayH8SrBH1sfy0wkfCkuwtw
kbOk7yJ45SOtyYcDVGHYcY0PhqU8sEcE/kbm4Jt2Jfb2M7bCk92RhoiRzxQtK99lViPy6so5aVDe
W0dn2cygK6NctpQv80YnykLAwPthGU+f0veAZezZjpBfLAKEIcSugtzaffFjoahVyvazQlH0IIHW
F+fKx5AsTo4ZE5SHlxMPurSwFBfZd6Jd/QcpR7OiOetLC1OgxWKjYSIS64OJMikZrcnr/JoZomIP
sVltjZWKDgK+2OCUBq8lSNPQ7Y4NgpsYh4DExbxC9JQgCXAkDsG3NpOxasfvScMDsYZlWJ+jmBG8
q4AVssJ+slQnnUMp346tV4EHqO2uxXdU4iscokzxS+yXy6uxWnR2Yjz4GSu9un/DaoXCqKtv5uuS
tEY1lsACgQIR7PMiTRazaqyTwuo7W/650Pea5CRtFxYYxhYiN9ziNMBBJKQiCrHG+zZV787pJJWL
wYPfQCXlw4p+jSpQnu6PzInRnmJf/LU1aTUgbjKTTWP/ZWAuKRg8B+J2LVx82HxptXjNzR2IEhoJ
XXRvJ3P7ky1UVfTmq2k3xZh7JcsDjxMLr5UVUxHotM00rY7MvBYHgTf2msmpA5hh9Q7Q9M/kGCwL
1e9EUq7ngjAlegXAOrFigt09aSx+L8GT7n6rnggs+4RhYEICfGcIoEe301AxFagp8yxiIGbzdoSw
IushM6UXc+/QYE1V1/JKHU1Q5q//YsCOWmNRAFu0qQgP81LOtaV1RlkEj55L+myk0krsaed+ryXk
dfHVoPgzqpqLMP2Dp4P2iRgF7CS+WNFVtUqNp5l7jEEuJ/1qQf1r/RtgDjSLEghBGhdJKOu4gurW
V9cX0/tKTR4ylI9VwDBTGc+C9DOD+7tCxY/WWiVtvhNsjveA6fg/3nYXid3TLC6Fa8dS33u5tWqG
5/8VoDnxMl7vMYG5LfN8Cz90EdovTjxB16SUybtosG+wd9ZmKrVqi2gt2e2H7+e/quuVJ09+vxFa
fDhuAwbU8ch3Kf0qreBh39Zy4B8XJM+SfNaJPNCdqOquCegxZy0T2v68YIlp8IUm2HAc01e5OAsD
d0zbmyOLc8XcNj8hWLxXDWHur7URJwVk9NhNxoYYE+b5tlUJZJPY8Q6aCbiSx7XQr52RflNYFDBX
FhzN047ehYkfh+4+feBhjfZ5VHs0i+VFdC4g8fKnTPY76t6q4t0fquwWUrGvEayjs2tCg3AZZ0X1
yYwhpH6xDrHiGoOzz3r+lRCUcgG3bJIIzxt7vZwSSjzbc/AejQrWZ0LtTgyTq9yCo+9YlIrx+wNj
TdbFZTmTzCGqJNCay0P9IxsbpNAaj1KWTqJrOQ+3NwyLnS4Ba1CpSXrkc6+oEkrbPFrDUljjn4c/
hab9LL782KFJzeA+7fcKQ4nEaxLXiJ+5HmjYVJwee2YL8TEFoKHhHSnwg2IlvVnoLjFmX4V+AA2W
wLN7Ygj8XHHnwmnfrMdu5A/GiTw313HUG29q3PKMbXkmFO0pawGgN9ZdjOiOWSWWAeE6GgivYBZt
fVwYunQS2GOLRpDzkipSS0sJ2+jxm6upe/ojxF6mtGT+sHK/KaPM2jvFtGBY7J5dWN5WKTntsaEj
ZM4DQQHyO7RLRw0m8zFKOOiHcI7ETSlmzRX/vZzRJDdb3H53DROUVFZR/ILc3OBsV8kwaWgzsxIc
8971FI3V0FfFazNISXRwPpUfVIueHKux9ecjJLdA9NVQE76El2smN4gAleNCjIoH06PJEnyUhM8w
0ZYSi0vtnI815CrYPrAAUW84oBh2w80ZbMBKhbGe+kFhF4gB6CQnUqo1XI3n71FrXzTNU0G8lViU
nuVX36vrQpj2sI+gK1Ifn+xHax/ZjPieQVYisJJ0HPLwC/CGUCYYqR/8Sedowh3LnkNb5L6ayEb5
4MwQcCMC+0LOd1mJzVqWEYFwlt7tnyDrRojKFjB5iC7JD7jyQeLd5JaWpsbvpiS6bwpkqX/Id35x
JYukaJCk1/a3YUwIP4ErdoxVUJPiUnUNuR+zlnTwCqaQ88InN9LIaX5ix23CrRvPMIQeDx7IJ8oM
0wzoNax+DSx5fI0pqlqElCNMx3ZgxKXNfqrWYZV3kABAP47axKEl64H6gKs+HAvW1/YjkFp5tWMh
xP5isdX+bwqRJGhWe7BqyYXkBv3f1vID5WHgY+fI5cKb4CFzxRwbkyq2C4jr0/RfV+DcfFkLQ3MA
LYE/mByB67Ucf9cOndYvStbi3cA/45NikO7V0fTLjQYQkIKKA4DidGiCpVvdGkY/2gurfPS5A85Z
VURUWZ/7Fshv3puTsKsKHGJra0wcCCID8a2C99G+J7eJvt3JpSCvd1PuIr2bqmaHpAFjja2/HqPV
YIBj6wy07skMmbDgzSLH3Zous8vMNcodKELFM31CrnJwm3buNvqEcQilyiA3BbbS/Iopgl6R/nRI
NBPkAEP4LSeuW0mf+ipauBZ+c7Mgpvmo46w0gpffTBjkvhL5+mrpY7D5zXTD+ffhvy6XspiaRBd0
SxpGa+qg0aeT+8+g8to34+P5i9dzju8gr28v5D+9UXux4dow7/dJkdZrjVHGDj+t98ktCqWuUX5p
IdnErbFtMs+dp45EocjStOWYt9LehhjkaSESeQpwJMmw3/l5OQ1kLGv8j+ZDuk7V4/5xr1vz9N8g
1neUE0KWsVmDun9NtQQw11JyBHWhHtBZxqu0a3w0TplXyBl2I64MyXucNt+iaCtFxtz045o7rpRQ
TrbRfN8mPmdn0fxL03Wd6wIJN8auwasF766OYPzisfeKQW2qEWG8XrYxl+eAUy7bAgBPxp2gx6Kx
IAW5MOZF1Ae0ort/K1CaRHDoV1DTahkzQnt16Daf8p1MTRwQrK9yg6QesMkV8Xk7tGBfSl9ipvVJ
Z+ljQhoPpKFx2y9CGq5AdiwHyyWJFXZrZ+40ZsMkNUpICbcHEvWvOIMiblWAA2C4PBq/CIR1+rR6
NwaNcaGKR82XZMG2qRF1TR/9zGsW4IvHj7VHhMep3JY6KuxOoFK36AEvWShK6dPFkkrGMNxuYr1Q
8BkBwCptA5omQEEmZd+grD/qu29DK3JC68AZE+MM8+a6dARqZ7AkDzNt/DfRmULANwuaiE7i3ls6
hub0enjKHcuiKx/7dVcyS91pdTwsBix3QwSfhP0dvvYpiYNmuM8TDtpdlTrYIm8NLk7Gnvx5o7tB
6lpX+8JtNOgdZofH77H28INgbJ6wHHZMaBFfOU7Si0DcFhd9N40jQ6gerjgOtxkktkfhiLACXR53
1Srm3RTUVOuhUPw9dyZL37QQSR+7KavNjetJKiPa1ZshyrqibMyexpNfjVl0iB+THcvA/VyH/ZxW
1uNuifkoWBbw2I+vwVQsXLrsgzCUS3KUL6ovtLYZH7EaqqcJuWFgJZZ46PSb7Lc5VkaRBsqPbGIu
GoRAH6gH7ym28uxBdhhWItpumoqBnB/pXBkViuAmRa8Jm0GFFdKDaZnra7u8TU26SjmKh0Zo63N9
Lcgf60UAtMjbY+fe/e5kMQF4MeBTvGKksRPibmm//PvRRRETk+nDfc7bBWl/vMCRzWsRt9BVNzwH
50eFtPLjYJtWcm2nFIqhCRlKhfHA2DNNqT822TbQs+V/GB98OQL8He2TYHkFTj/oSK4iLA0Xv/xo
tu35M4pHXJLvpQfKSMcXzK6JiBPIwxIXUnTTop4qTsLuGrBVkcpQKy/G1ovWPEV54syocHPcNGty
9JSF9CNFQLKbdN8iATgXozo3yr3iiifQqJ3pHvfR7sGRIZmRmsU6ATa7TxsYgYJHCzV+2R7GKcJA
HOViBTC4GykI/moOXj11OiOv2sjxqlljaF9rxw0UlztmDQca2vms2oFrt6KZHrbJVbQqOX6YlSaG
lX/vRdvCAWQoCQaunR5piUkbe6QOydc2vWklQHpuJjb4svBt88qK7xK0TeySjIXTGdtd+NQr10Bn
pKO/kfDuxi1ITIvSY8Qygz5pDbrITlYYNFTIFpOAfmTDQI3n9tSJt6NjgfIR7dVczl60em3FVboI
5fD2BfWv2MYnq0+3AswJejq6H68sJ6Q5nZKHhck0h7X4I5wjaCarH4sCTXYq1VhYTbxQugNfB9aT
hOC0+F8QydPUU4LA6kOzQkOXcdIg9Ef3/veNGD9SvBXCV+7R6Mpv7DsGFxDXH6uyJXKxTS4b6Uc5
L1FwSRP1FOsjNx468rrwPBJOQPJpNCfXvH00Q5ERbHkaWj8I8SLg7c1OaabZ0yd77p0r4V7vg8X/
PmFLfnHI5FHAIkfJefyztr/g/BbZ+ZH7689W37k8zJ+JmCHXv8CkkGm0YyMShmjcLFZycXcN9t6F
qSkNXZromxML6/kUqvgO7lU3V3ByNgXnRNh0FqgPK9wGD8aIxei+8/WgLrabhLeViy3RJtP+J7+v
jaCTZsYd79jg7gAiSAsvOFTdIgXJm5jWaMSM6PvCyzYwZmDDQgD6pP2iocIp8CWCugf6ka/UtAGy
Zw+VRbl/i9W9nwfFffzWUWUE0POB3ADrjTbHidCqichtULGqOMrq74wY3A4+tDieLuZoQvrzgVYu
jio3OCAhPv7OGPqXTdofnkZgHBsExwhqZpmKJMK9ZAOQdGjAPSLV2FrlokSUaH1LoF5gK6qMhEyJ
8umFCLDJY4msb3xSBIFD/65vzF9HrATHCBT9Fyd7VKejHtkN6EFYW69JJegNPqSBKjBuFPAeHwYj
6Gq9Y/VQ+80pZGu7REwUSkd5iKeXTcaP+QsK2n+m3mQaJkiwCtQm1iKdIwo95VL6hnmyFYZqgY9I
c96bRoId+OwMtjRb3JRuEhPAgLcT9hmHIFEP/K9Cmxy6N49DDoX27HCZ2vhNYmyPdOJ1t59xP3mB
gumwvecIXb0bsxaDWdX+5ceCUhnJGnOheIyMneuE6dR6ORu5LcrXbtTJRQPQSo6Nqr7a/cMMB8CW
8WZSuxr7ZzQRXxWTUKI3RDSNu3vLF8C1uFuKEQSpbKGLQUaN1aDlQ2M9OlaJgMGlk11o/nERDN3V
C/v8virTIO4DNXzNso00d1rvbkBCMtLjqsdZVjl8eDhKYc0/qLL+NLqFDcbyDEQGK5uf/iyy6dr1
RcpHaCs+EgT8CRKOY1uGy516rRXfoTZUbL00usUlpt1vFScWIFOeTyYBIhxLU4dw241lvBKyE/XR
wBH7XOL6qv+49noDvsJC1M5dJ+BR10DZa0Cgo+cGa7P1Th2IHnn0gyjmQEqWn/hPGAeJKemuS3PZ
YzdVxZuXHMxunvD4wu/6ODlG/Oh0rg0YNkPJkYllRL/feRREVhARTKujpPXMHRfZHNedK856jlYk
43U0J8Dr0ZlrGlN31Pxib69sqIg3EtwDLvuseH9kPrJ6h99/OL//0/43BHZmgLa6AcVpIXOrv0ve
gzNSuNZjC5rxAWWq8RuGt1yLeNL4Inye20ClHalKe7c9CwxIDIrSb8lq4V2PAoOsxiBN7e8ByMyP
kp9LGVviCjJhNDbJxWiIyJG0dpS25rOrbj0cVF4nOaJnzPIFAPTjXd7tjJ05770dauQGd6vqJh7I
awhN8ySQGBzYiQytQPtF3Pa850rzQK2k6cJILMq6oVsVrhIA3fPUR6falHfcIQzjMNNTszDkErRk
bsgvj0wTFO68JGnLFo0EdhZ+LY8J/sXSn0rtR60WeB46wdBp5jDC1Kd8HkT/N3vW1O0M9yz8D0IT
V8cRILiF7133GlvxMZ0YnMkogxlQA1Oh/+cfMW+TavjeZpIybC56WesVLbHI0gSBTvpbdthey1jY
jD3kOQJiUOTSSmtI/P/TiebnpI1H19/zBAqZMsk5RcvjM6OFTulYNJ12a6AS8Pw3Jt+BmibQEeRF
YImqxgslIGSDe41soGylqsgChDdv+9rbMdNF02dcVRQd1xYBe6AeasoHPWbIugBD/kRIB4lxWPir
wCqRxjtD+OS0pi9SC7B2X07rUcg+AKdUUuJIvvqOsLGLgyNv2+fVFS7U/WLLS+BmiIy7ntyE/7IM
Xasc8UQrEv36Wjbp48lZJr9upXOCxKsgfHjJ/HdzXVgxmKgpon7kTgU0NC3zLg3NSuJCH4hWYdCx
gPKAdX8weVV0MCnP5L0eaSQb0fBWoVciVsZGHqdekMzbH3ar5uB0lvgBu46n5XeJx4bL/91sLJ+g
lM4uvCXLb6ejyl5DtO2csB0LzfIOP3ueqmAvlvZbq4xolfIpSGNiMEGB41/bULxgP/UTO1njyZT+
YCOHzh1pKnnorIPzke6qiP/ytHI99zPTvyp+V8cxMxDDAz6jO7Fol50+WQsRSarrg637QM1LpuMI
D4VM5wAUnG5lG0zHpoheSlkEkaPdqSk7ygWyFulKVAufpogGYZmjTuiJlk8KFtvQIO8W8qxR59iw
3WpaImum6Qu+tsyWbYw6ag9RWQ5WXYl7rqiBTdaFRrGk1OClYXWRcZRbTmuaYVihZ2kSpH6eAEMp
CwgnMkwt6qYb9nYTxaOBEZ11nPYhuEmtcUfKOTFLj13KcoHr0CTYfmhMwO4i8C8/IObtfXUyH5RC
RsAZj2mIk/y2h4yM0OsiKC5AQiq5kXCmOmiVkFFzQjHr3y2j9L24veHP4WiSVhY8i2rljMtyhP0w
mmtVjkmqHAaDVZNR9egfKOptVBh2Lefbl0+Urjow3ZqpUFiZ6zg7XBl4fFOL5BuqDN/kFIMJUmIm
d/cj5rUpTXPx6j/tIqxw5pz8sL7Uc7T7/+jabAOq7GeRvhsDTrDpZ9qZn3e8oIiBln7a4JdjUCWF
GVSURVQpDYci5wFDe5XNv4mx4YZ40GIBouxypz4wFJklxhZuJnQveS4ibVGKI+9yk/TJxr5HVrQo
td+WPRdmo9pb9t0d69Ye502HFpUGbfriDfAk8lQmOjdURBKw5H85s9xnnBp6XuCghIPoOWSxisoS
jBO1jjAAIGalxamQ8Z9o8xQU5d/kMzgLdCjmo2OcknUWf9onrQpLWXqSYV5NpwHyVcWLatCFE8Lz
6CpBkvMxX3NPYQNyXKMe220FjzuvP6cjYdUN7WK8kH88Sgm9DQhG084hxqFD/kxzhZ/m4MlyGU2t
BU7ycdOEhFiJZClINEawb31IPPNdZ1y61jlyRHKjtf+0ySQBRnTawJMmxEMU6O3vF+s9b+LJGr3Y
RHDsPQj4D/6Wg9+Uo9FryPI4pVTc2clz+4Gqy4JNWhW9py6EQTV15AXBje3iY/8S7Cu0zhsRbKL+
/F3lLgedWza5ubVtJPiDcAfg0HI44UDGFvZClQ4tFpIlWW3E6Syh2DRGSnuKoIRLLDsDE6Q9aYWG
pdmpj1RWHYo1L/hJLd/BSMk/woskpTOO1G0uhF26Cmg2V7ZUEnbxdKblPAfpufp7hH811fdkccUP
u2I+BmVdkBxo21IUIahWQJcDlibloZMRwvRghY39NDBkI3Mo+UAVIhByfILugy7OD+yr15NyHEkj
kxXu4pphza2uKX/ZnbEjpv7sJomsqR+4AjvNq7kklm+0ttPgut6xGqtID8O4q6rjRtsdyHbcDyEJ
o9XXyr48zSCF/W6chXLguWYrxpavClfHYah5urq988euSs7wxtzhQpHkvMplokG/kCUvxO/suNfz
7BaaIh3zJNxpnp1QgQdIGwfZWGTEduXfGFuerRfDq1Hc+dqJlXn0/kl9k7k4tA0QMFHUEpdees2+
VkTEYhnUdzMTQN3J+szkoZXZzIIXMx3wvVICPs1v8pVwfGlWMmr15hddqgSnJGBusZyZyF1XTct6
FQQxSE1WHo1HI44Iiyu46kVHaLeTsjAg3mh9gxKx0d7H92+VnAegkwwmJOIQVOBhVam9bSVhvLxY
YOd/4IhC7qyzrBUfmED4T8yPxmhfyhMXQsEMPlo353LbUpJlViYPpeDzUu9EwYzmQ9m8FihWzD17
ocGuGApELhPAxHN+nj7wfwU2bOmXVZHPxWWk915KlSOc3ZbYykKIIapbRyXUMUMTPqfuROKCKTY8
D9ROyfZDvr5byrzTakC/Jowa6qAU3jpBu2DEiNQM2lMeZMibBQqf0eesHXF0SF6/dOoMDwL4Bfno
2ED9695tL5uQDD0hsEwOGqT1R5sVKNLloXN/kOrWbC81tzg42Dij5/8OjptxZgOVGqMUm4EXZgYU
vOk0nSNPu29yyDbYMN9th3UXzbOqeYYEf2Nj5DdFUz8PCwFD8IrS0Yq0HqVwmHkq3L/fprurR7Sb
upF3No6/tu6QPHk5eUX1UxiDqkeTiSsIHsxsZRoll+X39RZe+h9FWtiy85lmsPtIgIeEW9/l9Pbp
l3k8XUEbcJoICCZ8egslibqZQRmqipMpEyzbGv/V3ux8QlnKbEiuKYOF0m0TG2KosPbRzFR2mkXZ
34mw0zhRE6zTl4BWeXFHC+6M8cr7qkVOtWXRNmzHPt1g/BiSJAd/qtDQR2/8Q4s4W4T9lCBb9PuE
pXGCxOr/FmJ/+1cqyNJT8Ux1ImHNK654ask3KGChlL4WBaTqS+tMpYCptvhjBc299yADtWtf4OZb
lGjessm8rv/nFNXJPF64jleQoI6QWs0xyFY1nG/rtXFUyOY/zq+xK2kBhBwu6S7HTxqV2dIr+F09
/srpzr4PiiANu+sFmTq9YkEgHSCOxoZNNSg9QSdtyB20GQZfdRnzWu5I1Il9cztWKIxKLTyfh4M7
swkD9bTByXpb6fV6MAIoAPexlTgkGVWHuzfubR4o7Pm1l3x3Qo+VZQ3RmPkTf3DipGVpmRRju1ZF
my8hEfbkOmuZvMT5pR5DXNPvWA0CvHQKvckLLwoiUee5Z5K+mFBFhWOOsDErThX2dNeGGwlufKMj
Fnazl1/97kUvP4bzbW6MZQMQa/kcX4UC3T5WnvhzMjA4fFyXcCxX81pcyADv4FYEk15jY14ZJ+WT
J6kP4RKA4vvKHwisFgtvT/1Rt8YgaUh7XZHaMpHwc4WK9hQkNwiKgIIwlnHyP24VaHqTZBhZjrpa
L0fkqh1xe9Lugm8xpd8xMZJJck9NBkTsCKd2RuPYq4g4SgjPmBLdwJT+vERl7f8XIQ0SkkyjmP5k
QISLcu/inxk2ZW96ig4RoWZr0llERR4JEDib6RuUyzmZvlJhD/IEqw+xjG93ih34xQt8N79y//u6
8warAY/S2X4ZUeqS7ZXDqqOAjEp8k0zIW1/XLjwt0wYmn6DXbWrpfA3qM3YsLVniKRZP6cqTawsk
uqdrDg/WNyIw2VR2zIZJmYovPcVXJS/Z91QvRBMMfv8eDZG9kCJGpPiS84j71e6gBdFLJI5lsyUN
obNqNrNHHtYppZUiwMSw7itQ+hRwtKSZeoWLHXILrfZJd8CT6wZ1whacimp+6xuCqqmhglNekDmj
w3V/HGmmCbk0eem06gXiFj84ihGPgNMGmeEdGv3fU7TBC/ETmsZLttV/F0GTzfwEOwBGDat8Tg+E
RSq5fcVUcnA3fc22HJ1q2YYg2oIsPcmGOaEpoaTCdP3VDipVmbfxtw1+jrz0sLiL0vQdZBhjDyOH
eATNXatdk6EGE/8bvTRJ93h0zsHN2gpMFDPvpGz4X8jWGRHrO5ipVuwKFOkZOtga3+D2Uqa6vk7Y
g6nr3v5BtYoyqjrXr2OILOh8P6JybxVml+tmrQMbc3ckz58OcighqxjiuoM88E2x3Db0eFoaCsd5
bGW7rcCuP7xacA8c2ibJuQQf1zgJjBSt24f6FRjYkqfS8CleN7u4qc6e6KwzTBi3KYvlxtEAnNSq
PQt0Qpdsb2oC91hpCg4VkXYKmdZOEULLatcQDV4gYt3tgbJsq7KEyWtZRZm+nIJHwTAw1gZsWWkg
3Ag/+T5ZVkUFnu8/HR3Cpa6cvGAGEgJAapJgBwD/BIhI+U4BFS6Bft+9RXvj1/pVq98YOV2SdkJd
MKkiXcRpXWMWXpAIVL/UqXCM8AtAf23jVlDo4Q3yd0r5seVPNXw9OBvFH+4/Eadj3emGWFh6YjnH
AXTVKLrwqm+7UuFljPZlK6uJPAFoxe4sLmMR2tnX7XsXsJfsQXnGRtIagdZMYJG34nyPouFcCTTS
AHDuX1yDYb6gwDdJaa5yCHTUDdJnYrXcw1Q0OztdgKlH1rVIhICrniLd9V6NZCRmPsxAx1llpMMy
JEaWg+2vRj2cj6bDXb27PgeEh7g9RS1gt7AC2gtjc4GyIuW+z5B1vEpd1BbpPqNGmO774w+El3Jh
vxS2ICx6FfY7TSA0w4gVn0dkc4Mj9+CBSU6F7Dhoe2MRqCvC+SFbjjSGqXmWLWdvf+kP7MYgymAl
ajpXc8ze3+RtOxgidtk/REfSTBTyW1TQqJSVTBHMhr54SIDs7jV8jtq6I+P0Es72cg6HonahYaAG
UGrFCcUwKZX4nfINa4InmCjGEewEDNhRHoZ6NHSQgFgPhAYTTjS8NQblHT+ZVvxfboZuq/SZ9aeT
ZgwSd+IpTH8PF87t+UQQaTnQzsP83z2AIxMQ3BXjKTIRq4eIpESBB662cQebmREmpyhhST5wKppP
6/tQvq4BotHZptbHmdRVOSPBBXPqz78AL8avO9nxaH4Gkh7waHjTb9fws6D0+Eu+9UGOWXitbnv8
g/ICTekhpN86A2nSrAxBMVKgT6/rzKgzcpvrTMnClzyi4FKnd1NdNPmxgQVTJYndh6AfTb7T0Da7
b9mJRn6gk6mdcFam6lBQT2yZ4badVpXgMJftULLjdGPV2VGZxOSx5XcTFnQOzfathacmExvvRAmN
21ubXmaZw7E9Y1bBp3c34l8NRf5jOjjYvWS4VKGVAWM6mj8mCM1W8KPlVWpAidfuLgDYz3YrmmS3
drPEq2P18SjFjNyVEXXbwWgZUEg5N+Zo/z50yDRajXJH1kSi4C9yXV0KiPRTSdQWp4oQYAP7pyRF
UStHD19kHImB03SCwVdu2xofm9TKUbtYtJF5uI2egiRTKIT0YC98wW84S841s2d9h3JQuxSgg99b
X4EyO7OG2WGgrDJC5m+3GbmYXC7wIV+u19n/oe+h7v47AvPzx2mZRTG/zMRo3wWAon9c2jyiJhqV
Zt1EFVqx0OEbryRWfnuKGm2JbBPANYYbG+ZBco/ws/XqU2l6TBZksyvMMs8ld1MNua0WYSueuVbn
/iUgAgl46Vhrzhne/UfBUK4KCT1m430NpeJM9cYWVCqd5NT+hqnUCQZ+uq1B9Z8o4dIdyz6mhXKP
zvJiVBWI/hvNi/M52A2RT0PRkXsRkbKe/EblHSdjxcZMGmo2rIBA5bgJdHPAQxzk6Mmr+QhiaQAE
sf9BqNxTm+KFPGPk6ALge/o9Gsp8vyEBs8jULGt4fy/RXmewVeuv5L0d5ZLxdbYdtPkjrAmRoqnw
hf4ngD8qQzHR25XVLwsp31bEmPmQBtOefs2Y6MWOI0MFdVLZUoDMegjVxpN2c1oPIFBmAPOe+uGo
zKFJ3cMs9OApAd44hCYS9FvUOYc4HF1Ryvc9zoibQnqueBXe53jzui+HuYA+SdbCyWYGQ6zzrruW
/O0mv5AOsMeFFUBaHLgxyENdztnRTx3is3E4PEK6kHTiSz6OTmB1v8JkghDjTDCXP4ml2JnNfP/I
p11tj/NCn2iiQWoNWnUd2FLzCAZ7oTCgYK/JGFJcb+s5F5X9iaGVAVCbMcqdI9GEquWLU5TCVrqz
rqpZlYDvXJAuP1CMvMzBHF8uMR+fX0hjiZRyErLq/B+Y8KJuJDsDRKrwz88b8Jxn1lWgaRfxWuD3
rAtVmmSPdZGAzQFbqdPS67lpcCnLX69dbLMM/wUfsfYchVarR5RAJS9I7D2gClID5HmCnTpkXOl7
g/ZG4Imzvz+xFH2/H8PmIDu0BHTae1ka/5vhuBeCgdAco3EI+igXTZRZsOTbjjxN9BAO6unoVNpo
WWnNkl1IY9d0t+WdM+H+92FgXfX+J4DkqZyPHbuCXiG0wVo2NRDiZBxy49AqmEng7cmLMGQVkYkm
LpTy/YpRf0P6AbcSADWMoAEmj2+okVRmff0R7x44cccDOfVF0ixT0arxSwCx5QWNT6jt0gNMVAt7
4ZSqV4N4TPu1hpJd9j/xTbtIY8VG9ZkBlTXgE0L4bzBUcTPuRUuecKxrBJbuIU7aWiWi2qU3n605
n8aVvT56V05Dn2UkkIu63bIqYsR2ZxezJhn6cVO2fz4nM71dU1faQ6CwIPAjl4nD/SzTrYUZtvHH
Ul4+z2cThFWOqMPZ5UBt+ayDDZwYq6BiF6M8r1d1uwPl5NUqgqe0gtHJh36937N1L6Y1mCTISi4l
Ug+Oxr7W7CUiIDlB/gmJ8g6bH3GSCFGVegKLz/vbz9d+uQAEawyAMQTVASmohT4GV8z22Zbdtuzv
qcG08olOXOF6i+K0kfDo1YXDmmaeg/WQKdJt17Di/MRwKx+lKXVzYMoCqbXGyi2klAdOPqI/T8i0
hkVH4vHau4RR3F4EMYhxx0JKFfWrIGGCnC0LE/AOf2+2wfyHFKjg8qFK1NQ9wPZN77zDXbrkLwXG
7QiHgTA7QtDdNH9WTn6rikzlIMHK4oQ0m2kD5caow5bhgeGuO/RRowX+UcBr766xMRv6m4zuRFKC
OI8sHQ7g68t78rQc7tCqmfE7Y34mYlqmP6xVXo84eJZ4f+Dvq9qE1NHDRlNmNFp6Rv7HERAEZm2e
xI56pkQVMIH94vRdXu4LxTRaMLU8Xv61tgNYhP6e6X0KNL5m0FQ+iHJHdTF1QSQU8ll7QaenIYgQ
N9hzqpNyvaGKMDD4kQvVLm8fjMYpqg7bEjFkXTvpqIjPFajg2KLQvoXjP8yEcsZsYFH0wepqE8Wr
LrJz+IzBAy+E3bpQfkVr0UQkTZFIA3L8D39Ktfa3h38GbDqE6vhp5secNr9Z2gmIhdYHMqzLBFgU
Il4iCFABsnwKM9sSPSMUKxdAQczmL/k38drlnhJo0k/WU4gtvdai+CiwadYwdgFr3sAOp3iFPjNz
M2u1OSUtaj0x6hPsKkMD8HV2QAj+PWvm4+5MciGfPXnaLQjiRPoWDvsaC4aV7C5bxzZ9xj5i87jo
xSB4JzEDxzLPwjqk9Adlets0wPNb18xEF0YoMlT+VLKxi/Pl+AvbrzpqXl2vqiZ1NTzXxdCu7XOx
Fkx00wVlAjauI4sqeqTuBC5/QlTFnkyv0X8RSaAtWuBUrpJCPR0MsQdUX1YBsccH0QOwzDmYcGwb
o8xcPxfTSGgeqEUX/VApImKhNsj3wdvy0yHKhjU2k1DiX593OpKofTru96uolK3WHyoOvkX/OHpQ
QEQ8lDK7UFemnr00YXT8fhkAoqn7G0dp8Q+YhZa96VM7UvbtRV0fvxAhKrDzcl78bDGlT8KonGf7
mmHUemqlsfwYx3ljquMcTQfB+IjgGkFMgvJO+oOcl3HUExf8mnuBnTVyWfjMskL0n8aI3XLvfObY
I7DHy32hqBAp1xYO1CIwy/T5QgbFJvRKsPK2kKj1XqSKM1i7uSsptGsux/fjsMGmshS+Rwp9x47G
WOz/mXPeF1N49jFzaxpESR/o8BTZJXorTHRtcH+jpoeP7UnyEf9Ph5s4TbpUasJ6VT5k2iZE+zrB
X4kbOjqg7GS1EFe/UHXYmg1HhnaYse80OY5UTVyRCKcoDZtnQcVFehQEIgDJAcHfBb5UfWpaQEE1
fVRdYJRxC5knoNPFOp3iiLNm3WDIdYNDNUawOTH1fR3sM/y0qAvhbmyWiYbdS8xuWnd9obvIcsMK
JQAwVyJcKFucxbCFJ2IpbOpDkEKuh/B4q1BaVHo5iox6x4n4rty3g6GsJ9nFiaqklYLSCo0PfwCP
UZ8Nh6BO7L7KX/ybhPMMo0pxt2PylGw+cr1FUDewPT7uQRYD0wI0sWZhrOBrlp+ppiEnDcKgqBXA
OpzKvvoz7TL88kW5jfFbxEtgGPXHbXoQiz8Pr0Rxly3EiARk4EsVQvdbBn5Eaxcx4o2vjkXUPRpt
NSO02FwIwwN2vb4toWMXYQG0s0CI5Tn38r5qB9Vope/bSxw2Km/5+PBMdcbnYWkCpGe68WZWHprn
dvbgqPmmPHidT9vmSJwDZBS2gww+k4go9EotMtz/zd40MIo0ISUkTydTjib8dlOhh0S+TKNPqd+3
3SawNX1KR43hLjVLrbz+nFeeRvK9p4qdtqFzeVt3uB18nhtHt1dP7xJXAVN6t6lNr8TGMQAYQ56+
XoMnPTVD4//rMPjvBFQC2TDnXIj50OuTmKqcJbYwzZdJ5m4PIIjNkECAfc+Ip8ojZSFSggHOMzuF
U4MBE2QbGqAzJS6VzxuhDfEqrzHaj6mUErNZtsf8++XojxGDNFgPQvJus+E+HAANxQ3PGiAZJf//
qumt1BULx/8nVZxL0pKklRbq/9+DjChXXvKE0uUtGFO3MzwfuOiRHIPpkdLO5yI0HJt5cBsg1fXn
WFgraupqSRBTrLce+qgtsvfPHMJkc2xan/sSMJlHkqyluHkQzKJPkq2lgtRQk2AWXwi9i+fTBoaB
hdYC18YcBuZUY5sjVHh1ss6Fu2akJVlljUJnySibVVHjbPbNgugkQ1M0hQlRiocmDgl7L2Dig6K8
Gz7rqmZ6clNNIRZZaHzLBfRz2lqLQ4k1+r8l7L9tu4o5SsMkbxF0JUldGOjf+3Z066POMEjwdAxt
ygCrHpYmQ4gGXV4rwt39UZlOLkMMnp9V7MzZEmzCiy1153/2sTpBoe90TTgGoz01XdDVBwTAyH/p
3I6jxWinnMq+UFQb3iJbo1j3gLn8XEriJKtIKFv6s873IufF9XJqcKuT4PItK/eeO4zEpJ89lLS4
JE/enJiMbgSasXJUoq11T0Yp/2DGNrCSzdrdySPmvTNKOxG0+OArw6E06gwxiJmlbytQecm+/h7m
eBZkOTQULaQk9eZAoh2ONmEgvs9IdlFkNUqAXVTYN4rRPpNKaiYtVEa4WVJcyF8P2sQjDPC6+Kiy
CLKilJkoaR8bo1reomHoyUobTJiLEPBjKxrspsKkn3Z+PKVh+aey9s4jaRidZEdSgwrzcmtPZkix
iClOpJ5IV/N32Ah7SDmpj1V084lIjDlGHv79dvUbnc4YWuCm1xG4hxKm7XfvZMy/+7ejPry+cceZ
xxh8gRDiW2HE0NunCUAzZzdhEzZn/O4LUVsXI7JBHirjaHeaom7oo+NJGhb65f4ivhAlxukjUYic
jHux9cf5cwADG48Ue1lqep+6vRKuUR6BTlkH6h/iQcxtANRCOW423pIXQ8bZ2LmWMjq7vs8wCQqR
IMIf5BABOOghyieg5/ETZCMqVy4zrYwfhu1cKE+bdOMlT83prapCJ0YidSgvIN9PwxsTluMp+80H
jAcelu0mpksunofH96670WAfOL/Nfo4t4D+deFdkMQkb+FLuQdhymgXY2yLs5aISKqLOEzaPbOXx
V2O7+DCdkadlRPU5vpc0vPxIztJ5VnRY431m0j8R+kuOugzilmvN57ntZPYZpQlf24eFlzUVxPw7
Lduo6jjX7hN9aLzSFzy05YtZHblb7rdKBVGaR6u8QBwcm9MeEUjfd1BGv70NB8rCD8PmtMTbo/ug
V7efPDlM5YsQkCg8IeVlt+PpwBNpLEpWn7wQ97q6NVqB8krJdLQRFrt+RTa3aMKriKVdnO+cpAyk
Dnh91UL8yE8vb5RHRLZI2Ivwq0JYBJ7h7q/0kkSt25nrAjbswrQITZB7HhwExHUpilVykIcmmH2l
TqzY+sZIPj0YEu5iwISyVosamOf0D4vfvKbuDOzQ8gQrytQ8PWN1tW+PqguquzDhyUiWxBYIC1//
8ZqLqCJJRvz0nQkm5HtQ9pNvsvvgzI9OhgG3AdcisJmzyQEO4Ur9HdZjS1nbUBrfDl64spuCFSiJ
gZkKlutBrDo915wj5erQs6T4s74w3Mdi2b6YsILAYJGYl9LQ93169HQx1cuHNx105WSklKi6cPpg
Tn6LXMG2RpjUhgGkNQUUlZXiRdwvIUhg0Co43Vh65eCO6yAqu/N9d7jTcMl2tzKVwfuc4ZNabYqt
Zbr0rDzfYQLdbySZ3c+8g/uv2glYGvwYmUVh4XRLRa9TnQ7znumA8ijY1gKzL/nR1VvqsyUAfidS
QOv+7iB/aE70w5y2JBCw7QwlP/vcXJHIM1FiVqYIELFuzOx5K+hPD5bLnHJDB2gnlxGeanzf9+Ct
6P8vjN504AoQBUBmMksETj1UkbrhsAbrEjJrSFom+51L0+kBzNnXdup+Lb8e+2sdNQp+K97BHbW7
o8oQM0QQ1dqcN1ivugsqEZ7ntezxeuCcfzGAfW7P1/RNYyx9o8ovYyoDJovKdhFisxuEncSdilkJ
tqZTybdXh/58FbdvmzF5VutV/MVG15F5CdfiwKuM0bkqfI5TK8R2ZdcQgTI7vayW2r6EaJxQUvp8
WZWc0AiAXxNVPTVg6Z05CjOp+4cSh5ukx9ujMyOSUsXEWh+BUFoF803w61LyXhfP3Kfzd3WaCKbv
RPrZEuX6b2xS6EsWezpV2s2oPTM7YmS0XAh4hVksgbET0r2nIRu1GEBM9nX+msA2hkV7Vca/vYSD
EbLC2e0DXU4oY8wsGZrpwijc3Oa+INZKYHa437QiXO6v1jD2xg6LGGArOvvaW8gWlaZIb3W/W63C
TZX5pSpbAFqMhbOzYkOJc5O3vOPEx9b0grGUX9ybuvPxmSNyrTZzENnqCg0Woyqtn6D4+JzzlhBM
NnOZC3f6PW7CcR0qR4Sph5ayDQ/y3sghefFvoYcf86K1+yFmFFbCDFNjbjj5i95/Jonz7U0DSV9W
MZP2Oe8A4bhcm3Jkn3vTg0wrjLLCf6Kf/HIzc2wY2RwRVHIw1RrpY6ZYIpcUImONtbXQmXcvM/JU
LNTy/N8JvoWFUflwdze58/NSKydoAvBTtimDn/JKcA+7BiJJk+hv1gbgBgr7Bqk2MqxUfE+4+JJh
MGoX/PWhH8O4LINbir//MHU4ZGTbuj7hPBy1/2X9Am1/Dx8EdXR2KPgd6QWebR13Ogo3dI5MsOmq
7ghCgUpFtbsiqfYVudl/+i+B1HoXOB0JgdyD2UEwblcBcypEDezWFaXiX33KY2aRVgtuw99iyz3k
XWUcDVbc5ymA0QtK2RC4NnIPESQuncuwCaNiQey01284LDpmo1b/YGhoo20y5E7M3MGs1mDvxV3g
V7/9d9IHQZ8VRiP/9am/VKbC5w+ty4nqF0VtXgh/BwgLujBybDOTE4F+Xbc14sSEtpyfQqKyxi+x
KT0ADs1TJ5w7xhy5cvUedOkhsUELcGXXtzroGWwej5I6XhY34pFfevnR2xkF/OqayeMvSsPun4Y3
uODKOFQuErbMlWsn2d15rIzAnhCUO/x/BG7AUsLx4W8azorP9VfeubA6ZObY+RimMrTC12OUwIJD
81i8fxNYsIFvpKo3AH69Gm1jhHf9RhCLLTGHEA4TBj1ZtjrpwoJNiaisjvRM8fuuvHIG77zsGxAu
Xnugc/SKQwwlRZL7FFCZDpftqDTqgxDOSC2UUrBnB3nXDGlO7f17iOtok5I5hPSy7mW1e+W1alsn
p3MWytIyw5HiIHpsSYcMoyUY6HacX+52mJaxxOSUJtQA+oFmIsVhjHAgxkIFZW2k0+n5l7/2DmAn
JqvslMfbrk7EDd2Cpsr9T2oC1D4ws+2aGS4owdOSF18nqPktP4ccjyupp+olz38R92jGCuHtNpTy
GFe7H2yuPgStI6m6V+MAl7yWywpheC+VYj/J9aHZ22iKaCSXcYZ+7GpUOg8DDU8glAZWgOUgIQou
K+rJsKXzYhbpuvxHQ8Ovs65O22SmqqOVmYf2ZYRsW2Wea0ekiLdyb4mnL5Rag3IwIE/TVGawzJiP
mWEFYNXuVWuwMjLSHX20uRe6g5xrK29wTpFQvQ++IV5BotlcwVBSZFj/0CrNfTTbtGdk8P/C/2Kb
wrXoli6J6JLuIY+Bkj35GgjYUF3AIYcQ+shQhoU4IBZO9ztmWNdYMZNSGROrsGibZyhC7YxvWJ4x
A5aECDCgS4r0687nin8g6DieNDhmZxcNGYJGEw+LxzE2V7O8UP5PAcD9oRF4NzPGT+jgD+oJc44T
QolyefCXxiGt7K2lA4HinE4Shx3kCaJscvoEZumOfpQHTSuhPhemqWglTtLZZv1VZ13cBF8xRz2J
PEZ7sR/Iy/gAHo0s8nIMgt9GpadRa2kidun47THEzUezyi5hOam6waKYW6wQyiFm+Z8C8+LJX2fc
m5UnD58/WO7mQDU4UXTV+fHtvG3xGdWvsrnI8SQ/zyxyBqmfDXnnMBO7+opmGjIEQ95dyi8Is1Q1
hMsmUwmFVUhiAlINU+SxHDGDPmnA/wnC5YPcm/+xAYZdDvJUHOkG0pzlOkWkURalQ+B9++qQNMZQ
5cpPZEqtS432DmQO5zabc2gAms1p2/447u5eWw8njXT9HehTOeX74+iq2haReudjKVpoc6lOs9+M
+/qOufGo2ia9iYVT0INFO21GUqBHpR04rQMLwnJ3WGWJ5g5HC8xBdzm0bC9W34MsgvqgYbRMXYDC
WLSFOGp1pkQrJ2sSs5pOiGgbmPeBnv5s9rQeIE///dlAECFRLjehGp9T3XDUqmCtzbqZ2QfMFp/4
fpg0r2w5uGUMAxMi3ytV1VGny7oOBsYRHzYP2uL/h335UDAotx5P/x4Ls4w83h5fNcLzScs2UX0Z
MFeXmglxPMR3jgABY9FWaOBR57dGaoPy6THz5g1at965S1CdYo/BgWJAWZqfRydGSGTF9t2sbVOU
BvbTcbJk82rgN5VKebwUEO+K/wZMf84X3IjHO3ZkO052vnn8egll7FwqPAnYWY40cUAbeq/RMBkb
60yXNkkae7K61PElkNTsX2wHu3f4u/+XP4PvFuGv2tF0hlhmdkVnzXhA5GLUuds0NhfagHOHQ24/
++HPuubmkhehvYsWVaNOwQ8viNqik2WHWi2EXZpR8P1daLgFBqWzhi1IyO/xJLlTlWavbSlj4nNE
okJhkv5VwXhXuJGmqVQC3NlKirmZYc5wS+4Av0HDCAfe07Kln3eEe5M+Vmt3LeLjjHD0ZOxkIFbn
kuD+AO10UkQltsjaW81PYXO0eFJuY1/r2mt19n0kLe3E2hcFzsG0qNz1XCQowBhn9vH2+WeHjJc5
ieKvYJWlvo76DtK2ltB2+6oux+V9J7Re/eQ4055wTWod516JhDRPrXm1pICFltt+fcIGAtzRo7Mn
WmcdgeeLHVew8E5zVHFZ0pbbnM5mlQuRWxlVNbutgM/3YAAD745AioCUAyU43HGIaqGZrKb53XvM
BXQ7AP8CBBG2ZHF0sEGIqogUxF2Yr6rISjz/nH+FeFyeK8tWVsQUs+aM15iFaKA+XIeblNXfv+oI
SsY7MQc3z4arKKJXY18XSy1P0goq5t3A5E5qQ2QcK+dfWSgE0irRK+XjZmfkI7MshA80d77AD/gj
8ZQWUltNC+8uGrgsd/jv1LM9WETMhUL5I2xKYLRXxGDieuzcUWy73hqq6kQ5uBHh1kIe+hSSjwHU
HQ0bhSZ9EyEaxcIAWrv3OMFzQLkdcMvwzpQSr2zCQQPeqcQcpXeiN6IAsNaM3QpxKwOdq7uKlsI1
geUZwjZP4BxPObtM82s4xAzTZTTVeBn38DEkMoat1x1qWFuEIOi3pqvkaZJYke/7asc7tbcL6iCH
l6lGqrOkGjI9lnpYL7CzU5zLPPlYvIMcpRjZMus4rjibEpuHHRgYX8oZuUB5+5dEbBAuyTwvh9to
a3iIJtx/+APLArRcw6hNJsvRDQ1lPGms/JtJfVUDhYX1AUS6M1bpbc/JBo3Lwf8HBcMj5fF4crSo
PdccFZ7gng3MFaI8MfzrlbTguPgAuEuUXRT2R+Vj8lgiw1JVPeSbFTFAC7mBQw+3Y6z2RBXM9hCu
6SxvXLkFRuKPE6FZZK0xV2EH8Dt2WW8VER3Pi03FgLpoQvDRjVsXE2Nl/EGWEtmqBATkD8AxVygv
c9dkBw7tcdbYlUCeHG47MixTe9ezKc2tyOBNUDVuzbLCzUmuhCevi8EsPoSSzNhYmCME6EbwTfEr
xZ5dHF8bZVOn7ysdxGl+V96R4V5HL5LpfdsPjbXk/TIle9Y08oUU24JwbXCSRxaKIrdCwwmu6NbO
IAQVhH1OcUtBxab8B0mKg86nxXqTjCDZdYGAlN7DpL34Mt9Ag/UFGEpHBB5+/Veagrq7nuF3j/JL
jy3FdomEmFgjttilajU2ep4mqpu9b2j+NccgwmnT5rI4l2VSogdFrmlhOG/Q7I6dPcgS4k37v9yp
+g460TCcILIirxoP9w/FJ0O5LTh4rJYnu9aBy0m+QF5517HEDpQN4oW+htc1cTiXpWhmBMsqrMi9
ABFIHJVuTXHAxikk5fC4S4ka1IPPeqSXJosLjtQVgAGUKK6HyuH0tGqbqYHzxxD5NtWxg7vt+M7n
xMIouCX9TCEI9jiOt7xhYpmmPQSI/ARMelUWQLrMFEb2PH9+ullj+ZlD9iRRifRNbM9ozBTP3qP6
qW+2luetvqv1M3eizBJggHoDBAuFC6450xZWofY4AUxqvfBe7QWYMBxHrMSun4VaKVSNzbp3hF2A
qyW2/IXgeeW75rM7tUEZzvrNv8ggIn/4hOdm5s4Br3ANM+yXr3SBTX5SI3ckQM43e+NrrszEP+Rb
tUP6dVYoNzom8EItBF/fsCj4tbdovzmNUy5DYvS9nnK2Tj7C9xpkpLNRuQ/HYM6qZGAI4fGvxcSh
o5sxW53T+asPUIBY6TbDt/+/vddH2ZloRRIzIDxab1ikw9rSeTpna82flqE73MftbrdowmYdv3AI
ZMo/lqW2kkf6eHI0Vp11YPgqrfi4bMeR7NSr25C8MJmPJC5BsfiQuLCgKSWdrgZ9OJhgbDOiwJL9
sNqI4DIB0vc7UBZDuSiedcdIbjHwJm9IZjDsCA8CO1aQvNUmz3Z0M8qsEBELdDwh5pzBgVffEYjh
/diys3233uncIYqr0Ghu+PZkfh0EhIQH4jvUy1QT7KLVhnjxEPTr5ZgXamSaghbKoF2EjU7yw+aS
pDzP9ydC03CHZv9+RGWxyM/zw42hQbc6dPkZ+tOww347U2mhliEDHdGIY/O3/f4ITAnRq2FLdHZ/
OFKocrfl48WhUTZUxHAzeH3fiOgKbGP5IFcvEnu07U5mh3YVVv94R9Rrf5z3YmnOzWp8ygoCw0yP
1Hwszy5bG65jAUEzG3JilJc9wzB1FsjxRG/oLUWkA3S1HOzVFtwDf8K/lLBM1+R/wuz2Su6Qucks
PhwxSswE0tPcmMFyb7hbQgR7p+gTWa6twVXnX3n5piuoAENpm2tHbqjQ5I/2qARoB0PtqtyETJyg
PgbsKHzZs4Hm2IZqbBpJbjAu441OzW3ON9z/NBhqZsBkvW7NnivQXRnAp/1wXR2bbBT22HvGiu6k
yLRe7kq4hN+2p4HGc0lq6V6Ifw0rEEyLenziwPH0guyO0K6qzVNibRPUoiFuN642mc0mFkKPj0vu
Cp6+Zxv2yrLZ4uInCX4VEz+CJFtL85Wo1vvWhSOqeDvkcjcyMpGNCd/xXQutdLl1Fl66ff/vO/4d
LdFrXvAp/1CPacNzrolLLuX/Z2v7s0uwhDFW5n2Z8lKypfWJShvWvDqpX2J245fRte0vH6krv6eq
0og8KMgZ5dz1rohTD4lc5ejmWpDYiC39PDVZ5nTP8QeJugBTSgVol9F74pnnfsBz2SWIV73Q53LI
IsTzXuP4ET64OmSHR6C0JGtJRzWx2RlH2pTB6rBnNV0zmrzu8HWYwcVxX++hEwjTGEeyweigSidX
5gslV7F5BmvGbvUYTCxAyBsDRjZA7oVEEEUzyXWaidMSGGX/TZRJ1S9en+elnSGN7mrjrDuELDZ/
S5v5feprYVhLOhVH5DWtp83Jw3xPRyDP1/UjgSL6GxIJ2aYbiaM0Fwlkl079DvUBIdwLw826dQ5Q
AHEE5lqHAGZTHcn+iDxVlEn439Jf8I5b1BW2Uw2xYe1NFjMgRDzjwmnUUpj+wnESWUJba48eYLf0
3Gc2uSK+25+PioxWjLjpfJs4U/Fcv+dUINgzSvf6iNcNDgYbz0t5Pcbs7qMd4RovXEcInKAaHcnO
FPPzeVIeLHqwPB+TSaxUQoIygWCtxMVbEo0k3OzLw2QlVqN5VCCvQY423HiF3JGX4jAqKlEkvHUu
vdG1GbwtR0/r0VeAhLjV2XOz2J/kyLUCykLU/9fB8ef5SfwBhhcaA4/5B4wbhFJAq4m4lxUpK5Mt
cmZxeYeXP00fUPPRCq5lRtRwr/3XChyvlFiljFQJFNiZOJK1BN5ikRfZsLZU/rNFXbZ6U5WJ7aC1
WrLdtJ2LqLOwpwDX4py+2Wqglwe4CQdufoUIQLmARTVtlkvt+PNiNDIAMtFba3VXJ5kB7HrZ3SR8
JYcY2PPvfswf8VuGIJlJkA6AV8f3+qvZ3jH36lXXPTFZEmY4Tqlu7Jv/K5gDApdgSE9sdDj2hG1K
PZEIhqacx+ouR9TLR3bv+66RDBPOiowNIh2lDkGyBpVZgvCEemziBbkZTBuBUX46EHHbNmes+E49
DhvSvNaJGgO7MaI1chRynBeBgX8pMvcjDXk9+6wcpnFGYJVZv45nPc5rTZ38L54cXp1/a8O3w9u7
kw7zOjdsfX+Uqx8E3qD+4uga6nemKzYRDklVKbudNwqYBXNr5LiMCoiUOvzc/M1SKEAh1A9TLxug
SKERyJQJ23fpbhqzyELw0u2vsxhHYra2ukUqfjy563ggBrMtZhfP6Q+ro4pnsfRZMO5pnSzNB2Nt
rPt/RP/UWwMRF5Nx2h236LTojhKKGt3wr0DEWjjzNDOwMY7iUA3J/yOh6raLb3YE8+//lfChbMw8
BNi+YyQNV4Bw80OY14Tb/MEIXGwMdRhy1MhE/kGRAA5+768DS10M8af0mnNwe14sdGuoRTSPqhqY
FJ62V30aXrstJKMxJ0uLkUeA8iV7OUFLE2+NDtD6K+sFeEH0vriLt2E91eJOfuObB970bEG/sUbW
fJtryD3T3cMTHnzluubiEuRPjVLKTbu42vsIL1FJYsSoeQ7prnw0CRGECmxt7Z+u+IxLSSFRYAli
pr+8uETI+/4MNtzBc92iAdJ4KY0h0StDqIJPmDrEVboChorKega+ePQ5OJBGjB6ji4R2uF1ZCWd1
hmhJgVdH/byVmSTcPyUZbrT+hHTuQd5/vs4aWnlBZPC0IVRUuWfXDvUuu0I7dhzqZMbnDYyfNnlm
R7qmDuRpweJEBkRHJxQN6b8tyQW9rgDXZKpcGjneQ5BNUvkguCEBnlYyd7VaCE8lrQbkpzP8rBKa
5YaeDg3emv8w4U8sL7I3Yuyf9QPOtXikjdMrM2l5BiGjEsD/caAJRwRzEK3qpmq3qjVdoEXZidfR
ALQp5aUnCQa8fd9bdqcPlmlhkj9E9wnXzE8CQFruWnguV1nAvdKKErSUILT51vG7mSeho5H+oUq2
7gsP3xL6CKkN72oyQ0Bo8c7hTQOEd435HsraVFBDLOITP+Whw3aVzE5xYu0FgGJuCqs2vK1pocHf
FOFTuPKmJqzXdXVZSAbPT4RiDCy5zNglgP9jPtM4fjYHus0Kya0DV04MMVfnWcneNoMs19XMmkv5
P6ChzBQ6W4Vf34urpqzmFexSHAUU8tEEtWU+CRabjoTHUU1JrVFGG+DKzAKprU8r2/sLZdr5kMZe
nl6CQDxeXaPnX9xqzOye5GoZtvMT93acApQlonZMk+IineT3OYFRwUXDJ1BhegfiutX7dOxf1rHK
KI/tRVYhrq/mslyJ5dqmW+SJ/f5YB+Dmo2H7nkOeFCuNSt8TUt9Km1yU6Pxq07ZOjfzPxiIoMSPL
WgmmcO2iEwQ4pL/1usRtv/rF+PM/VtbMbA0ILxFq2H4v4WNoI5mOi3m7ZM4PUPSKmaN8/PdiqPpn
zWW2+bUV/BXjFEC6e6AiAtVMvAFnpKoP4iCVWL8LT32mB1uxifVHcSbtfB85vc90jGQGFIdMsrvf
118blfIzqHZddwcb0K06GIHCOE5JVPB6jfV/WFPHwOyidM/EnP4s2cDMqdcG7yKdkP9c8zix+52W
jjrgnLL6wBaenZIXNQpn9k6PmvMTLlBtRSFMVGihkbc8XM0ybyIuZEvQBXR9dA/QONc1sfuPyFmC
N3U9KaoFEe+paXdTFebED3AbiPPJBBuhdgrzY4Z5HOi7LwzY3U53cCAk430GDugu2AV0WfT2x2k6
1JZLf2tvH1+yOK4DaIbo9zeaQp2B42Oh4QugHQCOuzs5l1xw3hsR2afNkzTDTJxKovD49sQSOGIK
ox3l8Frfhn9+xslM2HQtB8he3++WSfFguH+9YFn17n5BqgxN1Pg66+cAKi4Zs8DCVok84lqqwBdS
0uBjYg4QnXkI1dcO8p9VYnTVuJsX6Gc1KPiMy438McKgzfdkqPPSrrssjEBYsX7zNmcvV7nJZH+s
JQ7xYhObjO+vLj8vrrV+hsATz/qadeJgW5y3ZjmzMcbGF3W8ZxHNG5BrwDcM3Auk3lGmae4KFBSH
iPwyHnWuergdIInA40VW5mLsB8mNFQg167Wy9SmFHVBK+ZHjibuoJEfxdK3bL8MYANkhDmhbRKeQ
pLQp0RbmfNRaiutAE+KtLqlnt7yOi/SU9tbtI7cAN2BWMqrAE5JkCLyJsTLZ4LJB/arNHA22NsV2
/S90q/j34biBO2MV6z/g6trhmFlKsE5vzAo/k3smOjZ8hcQr4BJZOnhxCXagFmDgoJ3+YJ1+2/xg
TtGoItk/LAasYHtP9bCR48cJHftndsbamWpNCmKhfaePVe3Q9KPz0jgDJTCUe3oaK41EsHwK95sc
onekULZyxWPKH9i8FYlVmeB3yrBOLW5PNJkVTI7hRV5TU09VpORWP5USesDrvMvECCUUb0b+o8Up
637gYgrxRycWF5npQLXqYmjFyw5dNewp3hU0ZwJDWA6AZtBqut/yoHS1Iwpc5Y0rgAlirFnnF26f
+Cu2ethz50bCKmKHaKCwqF6Ee44V6RYI3r81IdsQznBsSMcE5ChZuxUgqIQMoTdH+0vyeHuVmpjs
coRBLYEBJfvCtavz/AKHiBkNM2xeQAIpzn4pvh08cV76GJ1b8y30DUB0iQQ60LRQGpMU6/dhjaEh
9LQA0LWZXR17GsKlEGt5J8e0TQUnGXwliANIS93UjaEnIay8rupXWtyAHCWrPMu48lzgpiVtKiLw
KiZwKT9SXU56Pq9YVUnIyJo5sekyBGiBcdsJd10DDeMBZvflpYU/upmwxoYK7GUCfA63LBi43uqp
q5uOvXhL777cupoxb/tTt7S0SrwJVMfjek028tJpASD+D1tx2qbNMIafFYHJjaTXcltpfX1zY0Mv
UrA+gokSpUZJe3AT4E1Yz0rVajmwfq9RSlX15B8xNfy5K6yXvrb7W9Zq4+IhDHlv13uMgnFBt9BM
I0uQcS+dKuBTWsLEMOlbDUiVQyehVvPKisSDPEUVpg8plSY7TDPZv5RSQ64aMlW2EC7UJB3lDjSM
HOs3qSlUMTWWYZSI5pr6mAP/yGSDDc4/P5LQFW2QkyukgzD3Jj40h/Y9wJQ8NT2oZWJs/p45bDbo
oBRdfsVMjWuJkCBqI0flXZucyCE6w829ov3cL+ho4ZSlVU8mQhKDV/DCFN9zOS3ve1FgTlyYneLZ
thfhIZkEG1OfRgAOIDYPG4FPLA4jaxzoSF4kqf6lwcr+ZfJq6QgoRwbwditX5NAbOFamRBRDT7LC
Uag0fLSGNfItyWdBbC3zTAjJuULdy2pFiKbT7R5u7UAG7nv7I0BbXGv/v6SwPrfVbzNnQT9W4VBp
D2dOuRezxvFWu25y1PmiJ70F+UilPzJv2IuvPs38xz3zlv52eFnWZV/URek++vCCizkeKQfb2MVT
LtPZwu/zqtiubcf7LZvfNF0KcDeTsWpuOIoDQ1Uqc2OzWw1RCT0E/Dm1S8grHY7qyYS/Y4nA3+mo
dj7HsockzLTRIBpUnC4zoXn5qUsd+xl9TqqGEFQHXn7fX07VpohVEszk9RP5rp7fJ5JvKtlg7yaH
n46Mc39kKzPCTMdzq5DDcrD3h0KJh5zX2M86Pl/dZEEIMoet8hSOsZco8QG9+W5WqUNfxYiY4v8V
ZOLCz9AvcctR4ekc3rDdBbP2t7av7lGtE69uRs34X6af47ssSEfM7o2XqFbVXHjJonUai304o1TB
vC2RBlIeZ0wWJuLWspuZohMlDHrqNTMhjaUozJ3fQQTrixYuOCXNgvWO9beqzb6HOrTCq7gLRaTA
Yn5fnLpqexfhJyKJdRr5F2uVfeBgCnU+OQRMdMSeopNJlo0JJJFN+5ToE0OYhIpi4pzzkPpFCTeW
7kydga/3UghOKbWKpw6do9aPgCsBqbs8kWKIiR717cAQb8IW8E+Tw0EeOznVMrezApJoghgJm5rO
GczhnV4rNHeGktUsPO4YS5RaKuZyyaL5fsSidqRNos+ZEpu1pQ+Cy1O5hT3Sk2JGy9dFh15TUqcb
QmdwyDOVsC/frs3+TIYgF2mXM1UZE5/7Phdyh3c5GOZFTeoMvDtMpycM3ZXcqHSG55c7KZMadCqS
lVpo05dqdY0LQWFGe68Y0O756fuNM8eV3gtwOcHV2BBWcARYe4U0bO1SF3XnOCAiTdElOpptaQpd
u343wl7cYtjCYEdybp3s/6GkgtYg8BbyCWsTlEVXJ7J6wXBxDFOIU78Q8o4rhSZxORc/bgoryKQh
FQeH+pn6eB2It1XcPlzcRT9XEsE72cp2jZceCx/frsOzs557eagyG6qJpYn1EGhcQsDa+AH8bXcc
bVXAF27Sjh+ueznXKkTeRtCAcwov8aSgdH2Bet0s8tgFq5Fk5dhf3wMAasjpxw4GylMDogzrR10/
XZa8k6AJZY+hjbjIMCkHKUNMhDD6duqrmPOY1dOjr1FJnYUt7Pie+nhskoXfp0v/79S8KwZ8FPBp
MPJRnsLV5yZqVkmw3dWXM444fepnFN/BtsKX/KufP2f9ZOO7/AOovHopiZc9iZi1a7MMs3jjq+WV
ykHJus4byDuw91eM8648F6iLwelyKBUQFYFwRkVjZhsnFHRNvp2O08kfgCNVCgkWRR7l8usodrrK
eHagqgyjXiFHzsfOQYlrI6pvi9XVbiTiIIz3EvcPzz5Ig4ZtFk77CAprkdlhUJ0SZg5KGwj+9v2Q
PHYJngT11jU7q6y9U89Js3+Qk9YJ47WWkvB4HcU8YVBaTcmaKaeZX8JsU7mW+z6fVRkf4sX14s+D
JIKv1/FExYK2kJyU1gKT9q6AHq3W6jRE/toxYrszBTGo1h3qo5uRpmJ9SOXrv8wI+R+ODDS2oJRm
6g2L+wpnKBZvItVyX0/xaBwD/6KmxkUBHbMxfulFaQEoSD/9adTaRoX4PV1gJlQa52/CNA9uUAPM
7S3VG7e+6dcAdrTZEU+kfWhihZh3JbxR8H8zRg9je/Vbc6IbNYWqSKUj/uNPgNiRiuYN9FHDV2tC
LDxehPukJ9CDDYxUe45z6/asfAmQkPNryrZ0S76H8owV7v6o2KLU0YtX5hy3BBhtGv+XiY4MGAh9
siEZ9/vsfE9wqmcoyXbuHoEVtc3fHV0ko1wP/q2Gab90GIJZl+oq+zagQvn9zey4ljUYiFfUrlYx
/zAR1zIIQq6V74EOa/2i5ZR6kuj3WnL7LXpWjrBDUEvA1Fo0AGEhzWvAOx/nIlnpSVSAwJhnzC+m
PARSYV9CB8KOtvq/zDmtvoNZYJYEP2/FHKYHj6fIrCmpEu3AYKsEzuZqfwoQ0CfJwcm9Xd9zE94/
ddxfpmWLzB8WZzglTAKm/6ws1HX0CLCHgrAHVcyfSZoqD+bHBuS41NWjsRI7boACooPpkbR7zfLE
1QSMqoCulL03fcbBFk4+aKXnLunUkPHJA5apVW1Bsdg+glyxzgMerNZ1E8mZoLNNJZfWmfh3bxp7
lE1dRbzwzyMdHS81zi90kcv2pCWdhtP7yZcr6J+y9wM8caSMwJJWlVco9gvHxUR8sv3ltcicMnL0
moZ/N/LPwMLwZm7Bb078Xqxwax4wfrfxMy9pH5OqwekoD/ZHbtXbCmAyaBFrjKFupqYQKeOp9npp
1TadSH5HOx/J0giHVm/v4eBtEHYnumL20q/cLTRotVARck1Dfefg7LF7EaxqwMLHn06AJAlsTyy4
IQypltINXAxjH2AsnvfM8s/VJyhM7JkryRXIKiG9wmp/cWnuxwTRaoziPj8MvO9KpKbajh3/iqOf
/rYr106n6fA0fPMFqmEkqBoEi0WvVG+kRlYYYk9GFetIva2eNVlAL6pcgk2mSgih/koEeB+AIKyb
jognd8RuDX/6KdWf9C/nfs7bjfJgxq9sIQN3SWmbdTKMjdL23Cf4r8QWnnx3aDfC34TYDZbYG52W
qhd3nLkip4nPH2r4i27krjdtLsn4LtC9RCuiTJ8J/w6NvKEHMm+k9rxJBXkNbk28R8rEoMskK1am
/00nCDjsD2aIoLYLCTS9pVAiFh4E04N/myT3IC/xxAf4e8eyPH1NI3PSf7IRSKGkEuxqYoX05rp5
3yDO3r+8vQN2x9UCL0RVUj8ZWNUk/p/niAS5FC5O5Cq1bi7O2c/paFqVuh91pNRIQA9K8OIoBRbm
IgDOKRbaIoahDSOzP/ZbI6tiA5f/BtmQfxV+k+0U+Doi8uIdi5VTeLG947bl7HDathyB6ab/qI4J
iWRDPixKiv6KIP+QwONyCcV9vQe9fB9HSuL5iEIFCRRe/lZphq2PermmqN6R+Arq17X28EFKvMrH
JvCawT3xJlD531DJdRtGnxYymZMvAlMyn0rS2kSYhu1gdeeMWjxVL13iX+UiMDX4TBHh98/1hX2w
9nt3SM+BC4vZy+EsLp5kRaxIBnLZUX+NIOtudIKQb/nfXU4PnqwWm6LkHxdbmJazjpLBxNq31fQg
0dJjZ+jzQywe4PytMCTTbrxTNMmP9FHha9c/9fm/8gsFt7GZzBB9G7XdSdFvsz7v+RLiMTWI6POA
FROehNpI5WQHEQm0sdMNVBa8qc9ylu+RWNPkoblgzZXtXtWBOdz3wxeYjyq5LwHFY+fZmR6S8/wD
EePzwZjbW6Gwnx1dxc9D3c9Af4AYUkfWpoeiyX+VfOYiOQ3EU1XeMuqSVT5oYyXJPxuDx4yQXOrb
3RpgPXvKvfmgVfQMbbFtkm8/hVJ/f/IXwVjx11N6bW7fPBqq4bzO3EyQYlm99/oIEFt/i2+WkVil
4B1+ESSlHhTcmehoxD64yWZIMKOH0/RVl+vy4mwdXEVM6774FE6yXqw5XCqVO1OTwmmhTiwD1j8u
bVmo0SRzi8iMChq4kqzbnkB0Sp/b8I16qQREiR6QtVP9J7tW+mWwWLMfgsn65ZdUTTyc5sG7APHq
I14FvjzEDSaHWgXpyQohSKMep1E14vieG+oJGJBVtBjFXFT4nmKFOGuHzU850WNLghTAU2q4RCh6
Dlp362fMqY689gSBVHCkpKMTyJWF6MIVGIhJj4EWl/txi1OA1RdFm0Yd3lioS/aP/275ryqA34XO
mZzcXdnbSt8p/R6HSasLSbZqJzKGZZlFmyz+AcVw7WZknYv1EoISSl1FpSr0ryX2VouxsCOzC1E8
QIMEqrLOPVYZM4bmt4lI3bHHyXoeSLK7GHivt81/rVJTZddOTR7sCJlHGYLy/AWISVopjlz2LVTY
N0wjn1EoFSC/U6oY7LWmJHRAxFFurlBhWcJQPIHWqQv9NTATopTx98PIlaIzk9P8l8Yc+DQqIBmL
boGU3CmnrRMt//1w1Unh7CtNmTez7+swm/crjbQNgbwRLzrcgj3Zaked46pcqxQcr95YcdX/vGch
1f8sDNkw4uVt/1C4Yl/oN7qgN75ZKm0hAeGeiQd1WfTLFizo+nD/Bmdrh6uWsx7bw8ajUYnc1GIY
JewR79FgDGLipD99ajjZFuHOWCCk5eze9B2+ip3QNNDiQKsY+VoXXK6qzV5olKboSFGbqFXaUGNj
dd5V0AcyI1KwIvOQrf0rklAinxcjQan+EAnqN4+x7pAl5tL1tMFSDuIQYgfmlACl0y4DL8hMFWe9
zSN6CizL46/Bmx13ciTCABMbWJpk/SmzzTt6HmElYzLAUh7qeAMrQ83d+D2ct5cOKdq2COsXBtgW
H+9pBS5mCuG0aH7CbABb4SQkq9lMzX2sBStUTDg6gB/RLostiayg1byFy/jV6KsLwN/un+XNMBBE
HhFfxSDueVDUabGGbNqqz/SyHlrG6UfKJe9PzNftjNuHtRLw+61SKtaCEb8rUMvzFQ6TP94yA1Gd
LF11WnfkhZMtGzgcqjE6gCUX3Ybpf3CRLNlbG1X4ZX7moPBEzhi3zZ9GS1oQWQHqrzvTK4mk6VbU
NITQkhp/ogqfO4oQfaFsFrk872hr66imtA12HPT4XdOtJQtqJp24P3pOuw6enWkq5cNdTsDZZh8D
duLzy1jQe6m3g+CKqGrBK8g2fI7fs0+lx0uwCj/m4jyjIvSd0fPClTFOHgPA/pSScuFKOX4Wl4Hn
BTT3CAFNCsstFGZbRxqE1qG+SUq6qbos3qE4oco2WEtC05AFBzrLJZaCPMGnF/WJQxyFw10BOnPS
2rW/nfM5GpUV6iha7BDHHy3t/cXxSKOe9+kBNyQsDAdyD0x5mlMiY1RHtY3dF041nuFIhLTKTYc6
hqxH2OcZaU2FPPxsDkcOGRHAcEIJxNZhXl6ATzxIohY0yDIpXv5EKcYx93j5QjazhfHW7K0rF8dt
MIqEl6FGxeZSW3fOLpePrxt1S+7h6q6FvrZETKyfZjrefTGV+TR3FVc0n/Csk/AbVSOIvhdLJRVm
sBjtSR79Y+cQErB0Re7E7APwRVpAC9PVohMy5QSAKbHutP0IDNvYz7kL2OuisB2GIIzSNktYWvCT
O+1IVAZbtxTimcTULRFmFPQ0aL2TIe50dBRoxyHVaa6geW7ljlLupvT9SF4bpYVIXVaJcWY7+iK0
ZsOaLcgPX3CZ8Tco/e7nG0Tj5SXtycjqy06f5PX+OqkoVa1n43GjR67XE0rXlZlnbVLN6nG5eiqw
fDvp8h3MqThsKN139v5p5TkQLcm/E2NB4uLUTVTd9+p6Tf55OXk2n0khB2ATkRR7qt4b90C8qHFp
/A6MhC52X6XntDiA/AvfEjgyPEFnbTAKGiKxBrFo8TohcoqHmknrTdSrDaExJ2pnfgR6sO0/H1i1
QKcoqS8D2jOQn0kwsX2XX3BgFvONIzluDCi0vkYmo9fJ+3i/NqqNEo2hy7x3aBPouwroZfrQ8ujv
yLoHZ6wiLxUaN6XvDJyj/Y2deLISWBc+3g0O7LqP2UvowIRtCOOrfXM+AKI1FOOcTGGdf2m+9wXk
4UZNEtqdiHCqR12plG7tsCvYzGnFAgXyIK1n5sqEgXjo6fyulj5gB+SCze4YlC51W+jBmZZ1+Hl6
u0649eBwrmzkJkdWuT/7MvdKcU1Bkfnk1oneI98kQyaSpee34WFW2M6TWdbPiio8uazUXT2rz3oi
m2IkTdCDVSFLerOxpOHqGNAtbuZIauJ31QfoOPW5dCUMGo2c6XTEVxqdU1rMNHPRCgHM2gl25FbR
VPifeAmwDWivwixJdz87zqemVWHeGIb4KiJOitYIeUZwCVCoYTOoyw0fdATbpqm1OBn/s9o66n93
wSlv+Y4idsU41HzBmo68OFHdXKgItLdrV1xbXpw/nVOdL0bPeNhjMUQzh6DFwJEluqcYcggLo4MO
dgH7CQubGOSPNT1G32DzZaDKsUS7jTqU9IgYHP2weNo2n10YiDoe/O4KBfb2e0oXpZ2z7PIRpDjg
gl05A/hV+76c+ejAFuJd/Ci+F6at07GXsf5vHqny+/aVcflgqmkfIgdF1Yift1i83w/ghc5xAQpQ
aHU/9RlXoMkDyNkBsJskfANf26Q+gP3iiOuAlvv5uxJLJnqnkFAGOO8Axw64H1uyCMHEZC4ayFxI
V23xiTFnf0VBi7dmNjYyoQj3V+dubf4Q/Zc+iwY8LMstVEI4Rm6GHoMcVTtEcAF2Raioj/Pkda44
ezxqG0Pvf+eZXiqX5yhJCGjyGkUbTHG3BH5+J5R3jsQpx4x7K0a8QRwfvhTUeNlNq8q/Zev+awzu
+y9xrwTWwlg0vIPqIW1F1iJ0T8AluBeTQh+syImh2LpTOoZieHAK527xCOxhj7oR42MgFJdIImOK
epzfGgo/PDaDkkjZsynZ/gTxb4/Q6n3yi5YlV6uE5qt9h9WM9xOXJbjOBT9gZJVqoatCMDAovx/a
dZo/pbmL7xTNyi/LQ2BZozRw98CpF3bpSwByz46NzzGL5xjZYPWB/Twa9NHIEqpXs3rbcskDmGkP
UGhBJdQ5Te9jqi2+Sjq87CUTBKGFwxajyQF/f0lidOnOk614/Qj29nvWUuJS4yUBO0f4pADblIYq
u5E4nzpHjv/BcmOON5OWhueSuiHZdpHubPAOsqc2tpD1Al7vxo4gRJ07R/Uv7VIcc+lterwkM9db
1SzQ5DzuOfqXaMbl5Hyn0gcPvgAL+AmJuvzoRlKUblZaeHmopndp9q6CkR87E/DqqfnakDGM1c+i
cDi4de0HSPACidmXRbx8EQ42ej9ncxHKR0mOmibtvLvxk2HA+uZXpMyh/72Jr8F7RxTxXv91wftW
XBOPFNvsLMbqkm0/wMrN6Su5+b0uY9SntC11D+Y2gLJzOFLE4lbkpX7lHFeJw0bLO9Jfs61mgES0
2vw//owcyZfOtgJmg6dbP/q3LDaXlvG92rk7KmyRaVF+l+SFNlmLqfmj7VQtYuIe9sB82YajyD/c
58OGZO4BXrt2LOxxGFBjCztSvpvhpY1VHwjMpOp60q7R/DmaCB/5r7FhQPfDw1ebydqSKUIZxAQ8
beJXODS85W8iyd4efoFHj3r0ZXX9Ki9f8hX85hhU85tuYytmQwOhv9Gssqa4ishpxrnTULqTRrR2
XfW3oHg6oj32oWcbYuDyR1SgQnHDzNRaTtwzVBQW47bG7+kZXRBfQO7XbJ5k4m0xAUxfidHo/Hlt
JlUhCgNqY2TyxjCtYcJRAqGzFix1tux9kjmAr4bcVETNp1xGp3Ww18eBi0TgBfpokNs8jIsLANpQ
Zy/VUJIG2rrA6rqaGNqla4ax3TgTbBBwm/2I40I/ZaBX9qwiFSxWtGr5cCFOA805bLCzw0vzwunP
2pN42osxF+0HpFEX5dLvxfkFoDQEooQfxUD3nNG864q+JKcIJVbq3jWjp3PC5HnvfdvXMv0KBuNC
L4jU9aeAokE2sljnsJnsT4F/X2Mzx/tPvFx7vH12mUfsrEQW0YaytEvfUQ2T8cRUqNGqqpuVb4Fe
oLff5lkAQlv80mc7AZFWhmE/qDaXhQrITzdyRXkbhQMX7egPwNa/YVvj6h2PWIbprY11BZ/S0nNR
REY9V2C8DGK1UdapYEpGMdpQ7QI/qOpRv3IlGKdlCZsy6DOJxB8jpiiO9GFE6k3rwDa5eNK65sI2
da2NFJ2hY5WpyTLYYPVinPbUVIK1envqjEHTQTjBB7Y0npIhj3q7DftMnA0Sto+0V7BIUfDMbE4G
15j75Zd2gLbhEeYrv4BQRihiFD0jujaS4NA5bYOh50qzYvdHHc5sd9CPCYa/64aatE3lisvdwdOe
YnpHIz6wwOungNGIVRTK/9F7xd5rS7R16iycef8ErHqVYf9J6fV1Yfli8D0HOxzCf0ZYMGur86hl
DGSSaEyFfFvXxxtULkRD8OeUzphFv/xyvFslcCeQXe3n8O89H2YnXNrjlqrj7M18DQ7PwJtVB/o5
nbHF49PORyKb9lp1P9TZhtUpwwHFw2MZxF+/lUURsTcWya8wbFR6zF4RGZMcmhcroeLyTb/4YjBo
DhKxh3Q1thEYjGZEGLJH0JxJClBeaW0wzP2piXVB+BO3bx1xDZUQu/AmUAEVfCbN+HYtZdGfkyAv
1mIdO0Nini56OKQA91SkmQSxD9JvIE4PaGgazddQKKjMgWu6AR+hH9hU3+hIcv9q+KrfqTzZlkFZ
D593U/pfh0YV40GRGrprW4nMlxF46dUye6uzPN9Z191Ay5zBrZmyMovMAQDC/Edw3qK/zIl3hkq4
00zixEluVzwnolGjorN77Dy+A0QQI5eiS6Orh9ywGcg8QhnonmbHD2ZehMj0ahogHdeWwLKUFQyW
Qr4Uf0/conAzGGPfnBkgFWCK2sw/t+ZthCelv8rspcEFPh/Cbdc1KHWKe18wQVzwtalE8Un0uT8X
FC4c3IjUa3piW2lAeurHuDVzkf3YgYmZcWNung4j+omgj9nxJucOQ1eYQ2hCZ3bMoPytih9ieCKD
xmI87ARJYF/xTheACMwZQMDnFla7ynw9HsCxbR8iFlxvQKuHXdab20VAPnwEl9Vb0OXH/VDWnER8
om97mcAi37jqfRxlARuO3i84ihH3LpTULjYIs0f1gxhYOHAaM/9fwh8VAuzNHbP4Yux6Grh19ogW
q9aKo/ETV53n7KlQMQf8t/u4LrsweQraaLBI1PGDPdFG1m/ByTEnsgrDTFinVXEQ/lLWnLQKOORU
29ZFayRBHPr6OgleEoeVWQOk/Wl+obAvmmku4vKyEnHJ/RqNC4PhP7On542K0lMYtyIUfX6FfRY4
nfSNOcAOCZ0J4P11LaUlvkNFgoU0vIyT+jCNUArwxwNVhEcv7Fw/BipqA0XFE7g0bK9Gw1mvEj4J
PUCrTJFmSdZcHTPkQr5g20nqotL2SySqhWkMbq2jLEL2FFLQDHZ65DdGBZXkRgR/b8/laDKfWgbd
rc1IT0s5FwYcUL6ZloNH1ZjfAna3d3JqSLi8dmGMZXvIByUoWpqJk/a9i1prOGGUQ8ilDvnoCas6
LviT/yJQu/HaGIFDPzXqo3lskzvv99pKCzDGxi3V9cN0aJWMldqr1lee0PZAAg46uakN+bE/JtWg
UWIqkp/IFl3Xb/O/QCREzRvZFHRQCLUCmL9zNDm9NDSZZn9dy04hXghualRJXuyJ/NnX6XVP2Uad
BEvHnfpuhAFUaIVsUYfMGptzkLXo6FlyC7Xq5xrDlOxiEoFX3djFwWGKuxhZv565Al7CdGZZvAqh
cyUscLsRgb9D0UTS+RXhaYkWsc7K/JTiO/88ISYvgMiTNMtQbrJvzLq30PKAOV2gmozniBgFiO5F
T/IE6zG4w92GbP0QXGsVGlao+TVeZVb/0+qqq/xonPrQ9PRuscBb7QbFaBW6I1VY6g3u9RuoJG25
+KpQKpxIxSd5c5eX5OS7udABluFY8oAjxR80IkHIVvNS1nx+JRG0L7XXM6Jq+EmdGzgqo+OzYBCs
T0mx/y29yHdYM/UktoNOVfX1xgOhyiXYjwmzaJjXTR5t5HN4lzc43rv7nhWiFZFjS59XjlOIu3l7
mZ4N1HluHMUc0EGysueH3xHUZkjKytsVk2d0mCp7xOWoa7w1Rqt8mY2GApuiOOZB/GyA7Y1jxHuK
TD4hW0ZdAkPtDHDQHzJZDDRrlxoTQJpVopdUWAiQgD3BiNJlTXAmjBkHDqz1EEkKHOjc4DieWLuP
RVvkVNGmeAIhrxR+Li4Q54BPFvGnEwCr9OF2hzwiR5oIBWJF0Kbyx41MnbvwShOUCdQ3ix33o6CS
uYSGEFf6YqCxboUoR6tEY1s6NnUX5AdGQOcjO7qAGiNazscOnYXzA5Rp9pfI4hy5jMMoi3s5RuDV
m7z/UStkbxNafcpzBCVM7f9eN0RELDpF3CZ1DIEugkGc/is58n+v2Af5AHdi1Enn3SFxaR8ZVQO/
QBrhsjh3XIhDUY9ms3kn/oDpOrIZ7eCYD+0vT99u0NNheSfF06UD+yFM8si2UgP5QIAjbWGcNsis
SfVLGnjckxlXBUlxPR5H3RsgPcA7MJYAgvGgX5GbxIYKxz2pICNB9rHA+KBuIcTlPtGk/nj/Hgp1
p09MZzWFTpWjI8ufkE7XMlDRXppv+p+MN+4DsS5mSURy42rjgFYRwnJ39l3Cd9tY8jnL+s0TLdrw
ycpQyob0BSazjLZ0vOcdwe2enx07knXnSDPxwCdmUtgZ/RwVNhylYv3OkXQOLhO21W4KQ2y6ooRH
tQjaDwm4yZNhiiSZtF9tuIcoeEk1Mr8i3SwWXXzCK7NpTeUwgJNCRN2rgCPlhweI67zUxsT8gkzs
EGi1pMJnySgYFvlA2l6AxqEXr+PUARjaZBH14tp0ETQ9Zrh0pBnEwifyPYu+vpb8uDJTB2bDWxVX
KWLNFbvwVqzrJ2AJZIcDbNRgCJnOCwmOu23J9GWNSvTQhzLzEA9JgkPtTwO4hjfQvkhIoOYvpf9C
10KQCPo9+2HEzDXVTkHeriqW0zeaOUkhkY17FSdTOelY4u1R0BMKhPHw3fVKvCZuWGLBQs86sp5P
9PgnkqyYfG4LTmbN8dbgz81jt6Xjn3eB6kABjGXirYoBh3RVQZEyBqcfvtuUFMpD9mSKDr5zNRam
Y0ZKmNhWkdG8EoKKsGTy3FNNI9pPrFYCPkT4jGJ/kU5CZz8lPpQTtdafy9QwlOecqcxhQJ5ktx4P
M6JMuB7nRomMmOSb8BdTMgmW5xw2YpOiLZuXBoXmZiTeySQYHbkNVHZoVaoGnumljdfMzeHPmKOi
yiFCh2ETzwHsE1tdl+FWoPUkooTxpiZdT5aNc2g4KYiSgndd8gpt0ue0XdkxipUC+kncsIYxY6+L
3DGMhrgRdshoAnUmsmft0TjyqjrkaeQOeSJmCC+ovDUxeb6mEJRP35kgYXLhU6rj3/bRi+Ita4Wm
Mm1JpwMJa92i2VGlh47zWII6OLIe6HZZ/H3D8gm84zjv7JXH98ev+8EFFr7fYKp+/ozUTkWUjVlY
tIbduwuhSFwpOOYCwKhGMLNUApM+BdBwPcs+jVSU+DcadpPpqroIzowhtYzRbcKYHjK/1fYyljjw
/Wo0WqN/biVaXfCMvKzqdYuLoWcN7okcn8TFpqu0YDPkkaG8yZPOFpNKOivUlFMl58uIT2MIXhcB
/8gftDTQkSDfg56Pxp6O9ZKMtwsb2lSCEfBGxA0GtW08CiWEyGzWn8Fj07sdd/AdYSDM3cWrAXmw
L0ZalRSX4y/PQzksXqRzU/3uM2LIzMAm3KwLCPx8FF0txwim3LXkgKey0jNMCrvKZxD83mqCGSEX
ziBo/tGIi031c1Usq4ZFUmymIRYBGOzZHsHt8IAoakTLneBHkIMilfCIGiUWghCBx2i+uio8/r2D
LIENymU35uEwDHpLFO4bTmQFMQ5uUwHdTMCdkQWUuA9euhLH4EAefU4DLpXXfkjqg26T26wB5UID
Zngom+DqE2RiSUpN4sNOJCe6OKc0SKbhPhmRAaw9qlEdlfOM+CF+30nD6j0l61hqlVodHmHD/b8Q
/jJ3iGw1xZd8TopQbfwA1xiVf2AHWcc61iYwul7rrnJObd3tFKPa1l0UQJZseqeuvuZCw4I059M7
SFjhwpVLsSmOwQgh9Q6xjW3tG6wwwYnuWJftrgYPbyWZA7tXtHl6ZZU+7LDyEVT1UiQHaWRpWGx7
jGa4tW1Ipw2ETGEUsUrnm9p44xahKk9L7gGq6Bs3kME78XTe9LqB5Qm1u8oXw7HWXlYzK4MkR4sS
Uhq8vNPMdVV8qTILad7Kzzm8kFodKmisyur1lVdoxHaEne7vyx2UdXQiFh6VL4KzKXG5hWRsFslU
IEh6iLQ4GeQrwaZ3JnX0AKDs14ZGE8OzY8s7BHu8QXd2tJO4zJQ+37sFz0YW/PTm/KSF0QHjDH8O
rLa2793Wvt9Zvr2QgUON7kFfFt8RhC5AasO64Z/4wrGdsnwNgl5fDz3E7Evxy7WLY87yBtmgWiE0
hryFjPUYq7S0GLPyXNJc1mxx8vNo5gJArSYQjjFAW9EPNSpYHTVSGijOBOh3YPt4x3Bd8ccJWbKM
pajcp9aSKm7ENK/Ft1vyyjdhfeONeMN5QSOuD1nDl76Jh5ddLX2KpO3nL4DC/n/PKEoArwb8FvL3
dpUlLQAjbV3HWQh7aPLcmqCpgwJa4AyW9flI7UXF+oipbluyRJH+q1JbxUS9YHRTwnfDNxrplRNv
pAlDI3Z49Tq9y/7QTWJSXzY5/IDmkpvdjoj+2Xj4J+auWizVGXiZ//dJwcJ0tLPepz30SbhyIbHH
TMs3ow+cZDomd11pAEcZTM/eC58IzL+eHe0ADRO7d79r1PSs5Cj/svL6P7WufOejXeaN8xG6eDWm
BNOXkT6N9pv8HK1INRsVL2m+7GqD7e/BxoyUYOJUa4zU66IL/8HOzg3uoLT8hj6tN9nv784Emk5u
2enOiqlOK7XK8P1YSSg5pMgKbT5NQ5KSRvbupAe5k8iOat7VZcNia9ugXXoZIkdvsoQsrpqeVabW
xjLbyX1vrdZZDPB3tUDgenWHpywiyq6TOq9KsNVceIVqozgeH7fGYot6QFBtkYp3DmyRuEwBcnBO
lGg6sf3PRDOmyaVO0GgTkVok1z0kMVUT9ITkRWgYxJl4soJ5bnmoyzdQfmkycO/N/T32XpLrk4C2
UpxtGUJve17Mx8I3llRj5nY5IK4+Vc9ZDFYbTj7s6VNb4aJzKQCrynNDZddpb0mreIIdb2/KhL0w
Bg/bJhrVJK4GO4GbWzAzyYTMcNTU1yKiRnhBADyFHQugnfjDb6zJ9II4TDhGGrBFw7+5aDnoJtdA
9wdtn/xYcbWX9PwU+EgN9nmz2lMm16rSIvVYLgJmZ71zzmacrKnO6xXEGkEjbhi52ORYXuKM7A8p
nkll3yhb84RNLGapi1EVwSolxKeVFjZm5nuvhT7rNRp21FP7PgBpq86ShVrtPSt1VIwwYFYoeUo7
iTWdpwEOK5XZrI59SDKxRZnE96Sy4UPCrmuzqRYYKapwtxEhEuBzNuRsrISaTcrR9rMymnl0jU42
brKcZDoVPZ5lGxlE1J+oG40F+eOJCMskrDvBlLu93G98Pn4GqIdVl/a88k0nMXDNOWRLiSAHTP1f
tUNfphOTWjIuVYTMlg9ubzTnGa7PXKcpSBST22cfYaB2wk94/BaoiuCUj+XzuQQ0gxbQzMEU8heF
lb0AGedjISPMuucr45kMO8+USyQI4ihrhxiXCaKoZmObKn6jm+SH1ywtE94R4U07vIFfkIp5n8Gg
/Edh4leNDSpQHJNk1+kV3WuMVbEJvxMLapUxAt8LE9TRxKqnfL21fvArm/52k71D166sUWkeLKtr
3OJ9muLbLDeG0t1x/oE9haUH7o1hTOJ84eX8AiPZ3Qb3auirW3mE8JO5gFENr+AJdqRK7NHPYGkH
5xuVdvoccGkOpP/aNavwN6IQb2Y+edPgUbDffUUvHi9d9IHd25oxidOB4fEdrZPjvRKcoAvZTBDh
LNQYko/6BOyTaf7qZr0W4emZnurLm/KEBn4XEAb1XfMqP2UHDQa9jMCgUXDCww5+dof3fYt36VC5
mwmInn/8Ap2lBVOyp5Kp8DQMXvbdHOoyYOS/+aHW/HV2uZDoAesfwMCIgHdx1kX1egK/ZECFUYii
tmj7Zk8dBQ3BCTtF/6yezl8mYi7Wu+cUNzlaCCcvRCICP64WsHc2vwHA63a/HMiMawJA+ZFxXn6K
q0ljGAYSQElaPRn4x7/6Bi+iL9RDDABuTeNdpgPN3IFVmGis1gL07yA3IzCHfcvnoIjwCXa1iq0b
bvxvqXeY9bVk+TgEgsdawO99shyg9ZsgGOcyaA+fHI5qJmBk/opIJ1Yjk1EGZmADrbTO1eVdxWIu
dzLpqPpuw9EkDOMR3iFUd9srD64OBMyJwtJ6DTGOrBCv+CIFNLcxnc5DZn/W3Li9BBIUH9RjJP6N
lqV2NlC1aqHr0d5ExpRRX4b3ZQTHWbGPqKP1ZsgVmfpr/UM9RddyX7MmA/ZHiab4b/5PbNkM6ayp
aHvQLmhJxy36e1a5Kr+MOUqTcIaWoBxx/F8fgeU7POZUdpPE6robr8gsdFtjZqql7J/atmiFCZEK
9jHfAqsAYKQz+cXbja5lycYEMFrvfwopwshymFNbx9LrV9fEFpXUWknp0aR0KhZRZEWLwwNxWZ7a
1t+6Xy5sRoKV78lSqSLOT/iq9j06UaS2NQYuS2IKAZYR8EdinJr3DtxyVGQx5mm/uF2t7poOfIup
WpnmxYahEwK9rxx6joW07gJHob4N0XoMKabAnCRzZbbVM21ecsWAJgulyy6/UJ/YJ36noSQ09h3j
5E3Zm7jJuJaYTDRvLly5hxF+ZHlHuXoYcCmbdLEnazBEqI9yPFiWIE47PpzZTXM2815Bs8w9wW0M
RbwiJrDDgLMykxi/+tc5hzSD0RxTy9nPe0dasOA4thvQqP5I5u3WQ/tmCcPJqNq9MvnwiC41n3Oh
4zs2GMnwo+ryOJCxlWoviSw8vGUB3i4fw6lxNJ2F4X6Fx5JOQoO/Ir1AR4oqgs5oA7niDzIgB0V4
BoXdSJvQElbwT0x4e46gcJp0C3i1N/Joz3vk4q5rQ8FA0v9DRq5X7VEJ81HRnw2v94iButkHbIaG
cxSSk+Xmb0+ZGnG3XA6nCY/V4ubH7zaSswm2VgPWjzw/EBhuRCkjPJZ9gfs5t9hbc9/ElB33fgX3
aNVNQ3JhsWn42kvSz6n4a6zTZHsyMdxaJc4x+4RNAyQjxIQVVhwhZw9EUw+CjGxzFJyfN7/R6TiS
us0EnUcqxvgixLRW9djVOK9bNDrmhVhMt5TDz7+ReooverQ6yp5pytIW7TrkOUCyhnOL8Dg07aRb
XiRnPcKvzOHHFhJaKM0OnYYO00NXuKDP6/84pvvpC+pUClYKBnR3EPe3mW1ZgItMZpY3JcOU/kle
8PkINFutRNVlqLLWZO4SUQHaROeggvwl5YHkfQW4+/S9foK0cKRuZX4cbzrbiG2GFVGEbjfy91aV
eJ3WkKLq0BGodi4zs5CpWoAefRsf98azOc2WDCsSNeViNtn4heeUpkVD3D1a8shsE0xtDE7XBT1l
JcaJyv/DnIS5Jy+547bfbREn1O4zno8FXtiJ+Kik2pCQkZuZOdTVZNatyLaWli8aLgwwg69AqAaJ
6qBqZz3Gk8XP4UzKNUvNTMgX8rLvg5UV9TJxSAZiVzIKblxhEHxaLyGC6du4Wx04KGvc7Bmvspp6
XzJlRhNvILwHeOqI8RN1h8Lx0DKRp9TK1oCece2Uv3sQF22x/ZmBysTCUZi6psJdehbtMG2FOBI5
1r2aalccmg7KhyajKAeHA8stP3vvgxqT1ujq2CJ5hv7vcXxkPyEsrHRxDfJILY2bfaB/+1cNaQW2
r8BlfBynLJlVygjlCDAeW3a1nq4oGr7FxLzS/rirbg3q/ytP9G0XKj23SL8EzadfL1mjZv/+m1uN
PASLtYgIIOvRhybnHlAdgvjg9kvERvWJEXXjiukdMd0A0R0z9ORHr6kqzGgnh+qhp6qfbGD+BEWt
51A/Nx4j8wPV6xjZtcFr4zam1KxXFZAmILXaULx8D/BZ+rJIidCx9IVYXTqGWkkKVMtalx65FE2y
xaDU1yp/uiMaUQ5GfLE3R6o7+llb0lmr1P2b5aBeiXuaG/Ge20OZc0sA5745M5TRadqUs+TMO6ZN
Gv7vpVbb1U8eW2peuWr+08UbKFl+Vr1vfJ9Udt4GAdCN5mm8HCFFnOmzuxpkARGK830MNY2mUJ85
nzM3/X8gVdA6gx7idNLTBDRkqx3qkMBjGWPrldZaDMQfWtFHsGl1cgIDbS4sQFUrFWdhozXTsHst
W1mhkfXar4BxDP/SPphYnO4GZgrK4c7di0E6+ekvyZHGk7WWw+NMWCr/omRlid2EXkCAYVYwCDJg
C4sYfaPdM6E61Qiuawfx7bSuhpdWWZLkKjQo+Mxet0kMHVTaj8ZGJlQV9emU6f8lNHG/yB0a9jIC
q5fSJbdoowOc0CeCniHswBVo4zJpQQlGCikZl5tK77SEr8YWGdxjeXWpvXfTWzaiSGt1LlTohvR6
TUwYmBZ2xEpFJgI0pgy1N2X99VbMmJ0uCYklQ8cmmZHtL7GhaUm851KkBZA8cb/5g+ukA7gYls6X
iyTjH+BLp5vqMtdfGLbHR3B3GXbOd91NOzfJoESznKUabL0mRWwKwEgnaL6USuo1GaDwH6Y8Eo0K
2WmqY79t/wICEan17lVwHqlWJphVZ9R/ve2MwUU+jbROF6r/FbVPb1XMTb7gWmh8KPOtik6CzIrP
em6lpI1b3byTaKXYNrU6xD4o+XiuKEBCUEDv4Bs4s5B2oYdSQbTq/xoIzItVX/1dsBs7tOoG6RYr
nTk5OvtDd0e/95ikkZlcZQVxBMdnvXXpCZpWhgfjcOmnwdYw/9dVDHMLmQIl5P6axgJ/c0sjWNUn
qMzPi92QfLbeWfxQJKv23i9lTpab+zybiL+0WMOx8kk7WPOi/L2WJyUPBWqqKmJE6aYW6swUFY3g
ylKlS4dp4bSuJjyr9n3meDAHWqrLh5V/09XItze5gfCRw489f/5kUCdy5fyVPRuJe4GaEeXFbZAF
iMqnFPzr3MBbXGNzb0aBqEoqRIHpDjWeBVd0kRZpwwrYDl8MkY6LpSUFUClATFdJik8bJmTx0oGR
EPras9i/SYciZ/73VXSKEngAx7cvFcpi8awn+LFPfYGgP6lBuqqTiWEogcL4DclhoyU5rwNln+HL
1Q8RaKC9eKVxjJthYLdLh3zjT5suk+kiMNQcOTejAGJQ8mT1SFzHFooJa08YYnOttyV3VdEgaqmV
NxyVmf8fEkgx71upuOuhxKcVyq4aqLq1lJA25A//9m6KOC/DOW7NkYss8mecTlKAicphuSgzuqDs
E0elMMYy3s2+gRTo+GBAp5JH1Sn6e82f1+YskkSwE8NyhYkkNfLR+8q/6b6EuVcdh6m+leWiIqHW
pGbtJq9Q7uNUQbSUitYAkwVHiG18iaBdI4ycAd4irwOfhm5GUDT5emYAOTkkiUTN3izJcqEcz+oK
cbz/5XFU2OJEi16kVerSIpv5stQubib+Ba5dXxOmqdBQg9V9pC/nHJdNGx+bFhgvj6V805Afm8yQ
UqU56XTBXw7FAYJ9ECob4KYzkrUQohJaR///nwtImr+YWq38p7Sz2Bvd7k/bLSBCPZvJAN2jLLly
dxf/EW9oQfkOeQPTjqKwXQGFHUpoAkO4RNbaco6EVntLrXawpjuzHmdSNajwndxuv+5Zyr2SLoHy
baFAB7EuiV4CdVqNl14SFXUSHj7frU0ZGz3M7YJoNwEubl4dhwhOK6R7HicaGS1HbCdc0+IWkVSC
jvQnqw6kjxVmAuJES8NwXuA1cT9pvs5C1OlZGdYxFWsvn/xIuGayJssx6TSMne2hceMFg13DFFMf
ZXiSugaXjSxTcg/ESYWjqyyxACKxWgcxTenPc7E6o42udzYYesultdFI0ucV2N5xP/sWuH2NTaLc
lOgDcHR2fKpnjxpnBlyuXOgguoizrH27ZowoEEVOqVmz9vBrmIlrZT51xyEpIIJnxGl0LmpVybSR
/KyY9ieLOkKlKWKtmCgVMqFlPzhlbIXgDqvUT0qcWj5sL5lZPlXK6W7Xh1ZJEqa+t9iG7IbnQ9Fc
aMP0ONhC5CtO2vj44FYUf7FtdNBwEBU3tt1WTu0SwmRmr/MtzbghmuF46ErynUzm4jvC32HlH05A
PRdx8t8/I4AIcGoTwz4/dPdtazF0bKzL9Fe9Iodt27i3Xt3FB75K6fbtT7dyP0CtTeUGBvhT0sdz
EaoPYurzbGHiaBia1brvqwM1OXUrZJJEI7itfke6F0j8s0EnmHW08BRyNr4hVhUbsY0wjZj0aExE
MoB+C6qW8i5b6pgFDQKkxnhYLC898Azu5lBAxXwnt2HjhO7sUNrMRd4O5o2tF5ybG61GkLP39Y0f
x3qnBWQ5Mjw0yFTi9BF37jaIDUpBy8VzeuzlUMmNcp34iBp6CbZcwJ+2sfkVsRDsCqJKjcwvyVDh
8BX4n7D75LdVaBJbs4wm6jiXYixodD7xjMQeoAllgYY58ihXfcBJsTHCGXO5LswZz4u1isBShHL+
rc0+mi5x/B+p1dL1jKH24HNJApjshm2L0JYe8tK2zUY6SM7T/x8v7ZGwrllzmThwzxrlB0OPhkaC
V+p5mIhSX59H69GjsX8+dG67QMRv15usGxsQ6th4Bn2p9MeQMolTBGfjBWFlGIC3HuDAc1P5I9SC
jM7QuMvmh5eI6iJQEp+WN30LOJ66NH2FLKPDDRTtSTS+oOXtuC8C9GxmumnSciPFXmnzyulxMYcD
NluksQBJRBEz/ZjEST6BQmbKqnQ6jQytrEYcHCBZ1xf0Q3ICL/nKerWo8kuTS9mrpaWbOckgdERZ
qWQJjq48pvJ1LMQLDihmkWfJUN1diKwieQr/FMH3O8Unv9DddzbiHM+0akuMpDfNQ4XRpj/5JSK2
8Rom/IRePA8dzA8j4KuBd7UhO0ksuVrVu0Ksk88ErPpkCISJQXvzsFexeVox6P67cmED05tlyVZr
RwOZvnse5LuFfUtUdA4l9+PAh9DRiCRb7fIOzIB9UutmrkpNgT5yGmc4trN6un22VfZxlI28nCEy
LslOdz8kSBTOfO0VcFkErcGW7VxrUrYlR4EGtbYSmrNQaNjGCnzvq0svEjpxVVlqhqObOd5WJoxF
7o+B+T9Dr8ftctl4FjX6ukerFAUvWuShKTD8waRGtm4ICqAxF/6oOeO/4mI3IIQv+UCJK8Qamce1
APSpJW9ufHocGFxWuzWPL/4a6SJhcZFRSckdlAw7xQkrpLAJl61RnELiH4ac/8UVBvkLe+QqelUs
GDOH37wAsxHMaLgDfX2hOtk3vkIRez5LsRN7kUPoG2okyKZjRfhQ3X6PMXcpn7K6h10q1c0G3fTX
VYLBoCLgdOiWQHkwX7fLqsVqN7lDewxhkeVapDnH5Lkymc6k5JB4txA4rg/9oetgfxdxq/FS5FXc
n26UQZR4J3HSm3Qr3Sp/RJSaiv+qROpfB5u+sbKnPv0+v7YAHDZ9vUnvx6d8Q/x2UkFnk9Ta8pVV
s6Pq6xfbHRgMH76B6f4g+BJO9c0wMoKe1+JjYLIjfszsJ4t7WnRqqS/36zhZnOcPX2l1QxIdHEnh
OcUGsHTlJZaUf/seznFKDVjPFhNOTRMixD0NAIukRsUv9AYG8/Om5JWAqR2KqiY4W6tyqfzj4b5Z
UPBegxGBu3DJcFMpySLIPNEzvUyK5bc58ZNjn1WDDuCo1qX0eWygnrX6XWLxjFQpGHQCipCGWdOV
o3Dem5HlIlaAKbjwjWml4kqsbRQX9fznRS0twFcUQcbDN6lF0ldGEX30QyGKoe17HDeUl3f967IX
x5BDd/BhVtaJ1Qk4mUcQTnpvvQAdDQc8qH0jMcgzIP5QOEv3A5R2Kk4WiycBCoOY4K46E33FsmSE
6j34Fg+q9aumB/jnPkujqkN4xPF9uR1uLrRE0KpXAn4rYRIJ04gf0BvSlOKADtiC2DYI7CPWgmml
+h64oOmP4akyBjGRmutyxSU3oLfQ1I6VTm5xgw1VCoYGC4i7YFdY3TmJFNkz4JgDLZMbl0uOwFOn
2NSWU4BCf31ddjmcoa3HVcij4b92fDJi6fUp6d0gDNEW3/PMxTAOoklA5deLsooOxsJIs4WtvcMK
K6J0UOcPFf02cmXg76S1mqAgVxlrex70LfcYH1rXak75/uqxP5/AdlNKIjyad2CjwyTEil2PXQdq
P6hK3SpSoeOyRWmAOSn4uTEj0LXuO8WtvfH5t49qoudf4pJyo+EQ0hRHuulw0yK2GJLTtASezSqi
E/36e5EgndOLkY7t9dSVeZhNYI0xtFmYTd52XCvOywgcnj7gjAURdNQPbeArNLPxvxKByIeZHsfj
a1nfn2KLO+D0UtgpkHIuLYLTquilwpvr1kUzTfLfRIfg1HGoCK1Qi1cePexdcVDRDkc3goAYRkL8
rKAXI1hmrC2N3DHRCwuOTdUx/kCye//G4jWMa0dDDnKzwQtwjBY7s8WbXrPTiE9GOrSs/5Kol/it
ZZB5Qzl5Id4wWs6aohgxQfxv8z5A9NU5KSgY8Q+gMxiMdHzBTGdteFMMABw3gDFGByuQ9SMLPmZr
pQf94MOGXhoBW/zQ3VL7BbHu3JgUMTDvWJwurNtHzzTFxpsAQRuqSI98hu08eYoELMI4XxFMNzzo
+WeDnMusR0+BF67vcTNt4K8C1T0kuIZSRMErHVZHkaQcQUUlCves8y3kyTXjSYUxryQuczwwfoYO
q0cwbxW4genGp1lZ7Kfabn6VH13n6oHyIFMqCd4V1LrsgduqRTvd8LIRjmdXeCaUiLj8UkYWwF2y
iHFT5i9f4TbYrzH9ToZJPctFp81qm562pjYYiy3zJNOrjXmN5tYhhdXCbO6jnYeklBXVspT+q551
1yIPv3RJzRLB/qBBvUx/eO7KFPz+vbB30i5gN7RfpxUzwPKSHppB5n3oEhoqRuIT/X2DS3faH6VN
UsmN8W2h8OOBOaGT3qOzhobPRBlqJHEQO8U/zjvcsi7ktelRDbuma9EMGCh6QdQEbiq9RjoQTJYP
96jNU07FpH6Idg551nTm6bjEyL4Gp3WCEisRjHrFxGD+ITxW29lnn5tMcA0quLwtC1zNzpCunDGD
8y7xyHmdL9C8kuR3OvJS5zaT9hr9DzP34HaXNl5f81zt5avRiStUzzf/O3xmuF3+9FxkKin1PA6C
tS/CZUm28oIl31M7xfS2yMS/cqc8AyXvkd/HdIi2+2p9WiKlx7WdN1AupeLFJnGp3Ve6CGaZRACF
noynCuW7ClEsdetXhbM56C6uFNY5uNyrFaMs2yHUH6WVXaf6NYxlCd8sMMo81aL6LqNgudrDkw1F
A9WkQjB1d7Zq/MCjCzmsJjudrJqxKKPODLMfnmoMzO1xeHi0Toyv+kEmoxQGuRtrFDGRfYuPjm1l
ixqJPDRO86ZxjFgXlFO/r7N8e/wgbTY3RAR6lObrVPzq7yKfIHSBkw72pzu21ZeC1bjAQi5fB3oN
9/VFMxn5c+EnRT9iHbaDAwnFpzhiseFXBKJYKQR2L4rITYaVxv4+6698qf3tVKVBDiUeDrBJ7VKC
9I6SKys5zNiI4iX4IdHodNT4zDujnOIBw1Tr8OMlnnSCRP174Yh7OM1k+XmvAAIFvBnRo/tDGlCP
sWsyDBgokq0aCLi52oBFGHzu6n/vxWU4hM5VPxDsVc4yRMufZ4jVDWDXA/f2h7AS1lu6E7Dg6xgl
5Re0umADzPfB+upcOXuyln8tClxgHDXacAnXtJjcZG3gbu0Hcr9hLQ3I8tKOKSVo9LA3RU9eIbTV
4WX4U+/pLu6g/2nQUojR9cdBJP8+3K/2BL5nE4EMmoH5ndqHSanwOxo7WPey5NMtXTeqqHvZbdz7
F+oJKCatkaVuvBWIIlfNGOQw8xVfUMp7fPmGURG65gDWb2GroGeowVGNjthf/4un+AjGK/QoHBc3
0gPgypJ/zShc5ACdUUuBIHXXAy3/QEDZ1GFYZNr2ZURNrkj5zaYBQYlfne3MD5qwr9iLIiY03qBF
mSBSn2s3jFdYRbqOyk5EqZw08SymDbASH2GJ1NsyZ3UHhXzSrMvauq7nb9SBTY+YLbLZeL7scG5H
PWbdWaZsz+t0DCyRteN/dtRvH94DdjwvmXJJLOefLzBWPJTES2ffYvb1corjql/muyymrFN3Y/gA
cFPqYsIO6R/vjl92Hp8Dg5KIR4S6mG4a0jZ1+9AbRlYFq84gK7ebOey5vjqVTop13D+V6JKFuq8e
s8i/W61bA0jKeo7kWEsB6vJQYSBAwJcHJmp3YsRmz+9oZkPMxYGN0IyOkMro3PyfWSM0zESbkjMo
JKRXgBZEyfCEnsbXvPaJ7X2/E7+TWxDw5aHPslyb7si++rsUJt7OiukLMisV8R91ANVpGsL+/Dyw
Ri3RfXk+hKbCVZ0U1kgX2liyYXdaWqnyv/t+qkyhqCVld5wzRF5CT+xlL7nd5qw3SKP9Q5ZI4hwe
u0H7W1/qKE7gbvlvcdOfsTHTUzJjJ3dnj7vN3f2CCxav+Hn6mKcxoJMBU8NFclEdZvsqSHWXOIGI
C3sVWTjFCvJATU3MEVT0uBVehS95vTpRIcPY6P39WdNtkUfRftrl+qPwqGxFjL1ftmg0+nsbFAHJ
+kEibyM+BCyFWCVC4ztrZuAuEnlLHH9IOMPMt/FmTtMZD+7EiRopD7b53i/xvO7jF0cPV24ox5Yh
InkDoD4j/Ke4G7d2ImjhFzHsvABmuArSpkebva0otJDj8Px+QYlBzBkLhsIO5l/SCzzSQI2kOM1/
Y76TLxYyMP3s+IWBYydcCrwn+VF+/2MzyTmkT9uuYwFC7B/svKm7xnUBDMWXtydNCMxCzAdQErXz
8NpJ3GN8mtGmv+vc881+WWC03EBEvz5IYM1X8d+WPrVSiTACELekr94vQ7YaV4AM30UlNN/C9FSn
efc4mBZ3Do9/SJ7yrybdikGm0Y3Y33Sn/vVmlR/37yvlHDPVG//Lc/1veFcJ5VwuPFphtyHTNUlD
cDMYbNSbkHIwGpTg9OE/dUXLdk3x9jaSQOx3ieo6F6xgAq4o6XF62HYFxEBP3jd4Y4IG25MYfugO
zl/EjWZ+1MmEknOecK3uYExpmLhcPM1HLewGAbp0RK6nIPjuxpCdBPT7/6wbhGpeHZcNZQYdtj+z
BuGecGfR7gHEE4PAjAZ5BfiJdJmONkK24RU2lMzEmy8mzHE0nERSuqDtyhLg5cVx/qm/bLQyH0+C
ATd0n68Qd59KOgQcGohujfX1YnlioNTJcez+/Nu/XzbbAXXIfMhkYbXOOz3OD4KrWKU585eQTW4z
XXg4QXKF4QCfWKlyfUcvHF73qvpW1yl9O5UfVcteV1NKaRNTskp5SPyyyd+bcj5jCBh80QJXN/5a
FwEX4TZWKwDFeAAlaLS0st/d1uJmTb5JVKL3Ow7PQJGpckxN9ahigprGafEP1IayyDayUcpxtc0i
pzOCJmFKVHmvRkF0zcM8NPpvGhH8F1gLudb2TTYhe8pVD/re8a+UU2CkmUZgfca2IPc6P9uRtqR6
t5/DFEIyRyxDis4ZSiS5HTjisOOcuoaX7tNYsuZZ5EOZoERqf8+VtKOSLP3fs8WpJeIH9ToSMED+
F6H7Nfc46ZygnFW9Pm7zq4bEYa6X5/iyrGqjQ1NRTHaPSsq6QnLZBQQSG+xjgMoGThThnd5bomvZ
E8s8koZ7ohCqeNuD14A6gHO2VuYTost85YXsfiGcmt+biGXpo+W76lcadcLGPBCf6E38Jz3mWKn6
biT3QL95dcNM9ie1GuMiDRKbeMF9LkCD9rEVQWxk7WeYQXijh04o8ZCOva4dymKUpSph/4RXdMgO
KcsmaPv+9fVLb37o82Vof8+WxBEZrIiNOaptRUGE+IzVKxsH5qdsXvtLZyOTA1NQJhmTqijfUEec
B1ftvMRROZj1O/+BjszaA97krb3R3tWGfz6it7EZ+N0CL9fY/3bWF+fSKHbEbI86t2HHDZ5KCT2E
VO3RcbrOmhjM1Zc+AYb2ANHhS1q8GMEZlZCMuM6r+XAoxrCfw8ADCbULaaHuVuhXgRiwUIUyKdy/
gzWq7GcYHUBTw6X7XyAipNBAMuR3iGpqaq6OJ1ioB7CKDgNdCS/MCR4W2TwaomV3DNysye+EBwnS
gCpGj/kH0dJPZvuFxCdcjo8D5d0Z/bw89Id+ivFHOaYi66w8hk4wHxwZDFYQg9LOeB3kUk30wc/d
p9h4eqDEfnyJVHjZ8LPSdgp3HPS9gGvPfzVe/OnkCdGKHSWll/hOoue5QCscQljcRyAaFWEHt/0P
WaKdOww73vuC5mcK9+dDTyxZKGXWXPSe06r489UyQlLN1t5iyF7wKfmBWI+UCUSRHQ/0Dis63deP
SqKUk158bRFmp1/kDAw8aGbLOJ/kbXaXr3VtC+A1YDYF9+NOe7aDViaqBT4aGADFPCTafcGT/WyY
RqwylVNsuI4MgQCb1uEWMbgqqKXmC6sF7Ecinkw7tPpCLYen9XvTT1kz6BR/+Y+xuhWVxT0fO6Nh
FC6KTHxQLIJSi3Ml0oZbR5GusG8tKySyz3hn4vrnVla8I91E/KW142VYaTtLqxbzulKScFGVC2bu
E3A2qF2pJln5fyn6kZ112zTtRqhrxfG1K8ucjzANkrpLKQ1bahweRk+gvEDk/Xo6vw++6zmbNKvc
L4lPZYcAb8fFLCFDkJFeVMv4ADA6z2cwlAmGsXNaIZ9la0/rD/SULW/GoglDQbDq0NucxqoZZb2H
nwH02ZcbeIz3h53I7YmBOO7rn2gBRWl0PWkMIn2X/pKmJ1EyU8c27W4QNGqf32uYl/okKTA0DIaP
gTsbbfj6rV6sbVaJUtEVYgFf+lw3zBmUcQscft0r/KrEGzFPcNMKFk4z6ZCvaLQze9JRyNXnTlCm
DN8gwtBYUz6yCyVT7BiRqfnmeaXJ21WfHHWl5Djc8KM8iqQ5/X2xVI+5e2x1JXcFA436HxwrNdPA
0mi3hXQ4tBciclX5y9GD/KdrN39vpDsq/fvfLG4hwvRUSEemvPSB9VlIkIn+2ixQkPxPaNSlkXJ7
XScIQqQz8lRFkkDkJqZgKsK149lP3hhqjjEBWe2U9qy1DeQ5M1jfv8N7hA6JV8IlsLWt6FXjWxDu
vc+zW/USb6gpoQSvMKQTrE3DRLn/MsTY3VLxh+h9E/z2NpSvAvHFjdHBFIE/GgG9+gA+xvadbckm
2Dd59xbtBdv4ZihFhTP7knSc7jZvzhxiG4H78bNKlUvbjZH5+atUEMbEnpKhkX11aoriIkt3yJpW
6/ofMgLKWvzFow8kZW8d5WX4uV1LjsywAXp8Qj/pPOnIJ3p3ZVvK7+9WxIgPJeu5rkE6fMGhmYdc
EsssXiBZWu+zgYWUled7BZjVrExHRaAouZ67vli4PcYSqJ06m4gR7S8zieMkY+bY/Lv5R1b6DMue
/SV6vcVKrEoSjXbHyNg6KyI0CAvsspE+4J80ARAOa0cNiPIfC0hrtFbK3jBixlOFf4fSak/5XMjM
rO3G6dFXi/1JvR+Y5MKYDeQ06ROQI+i+KmGekInxHLh3ww6j2Dax3KUcNngySBfzgVkrhJ/pl5D/
osiJnOd1Qal8k+wNC2a8fSbKUGEaeDTpAgkCYmFg3OiJdOX3ev7kWPRRo3w15TshjegUgicAEE7+
GOUZC0XbITN7WBtOV0antVYgHen4aFDwrfHbwoAoiP5VeH/C/mblL/1W3Fwrk+9JTE8t+qGQYhzr
49tdMzViXQ+Y+DfWjk7xF/S5Z+A1HU6auhLoBk8bozfSRvZNOiuwMTi5MIMxqINBRIEwMEKmcLlt
eq7OBEBJ/Yn5uzkh2BQEfzrHpLHt6p+HQGPqdtBwhLsaAuUUz4jWSJ93NGFxVPWdPH9TJQdzBy+9
Z6xDRPH5Krj8du5DSuYuf+oQq5PZuwCiqqM0gDF9FD0eoOaE8nb9Ugl8BWrDyLZ4AEHx1ZruRjgD
R6KyohTqqE0akrzOkON2qzjOx5tcZPL7ja1kH602gaUYkZlWSsVBX7+SrGijibKPipTnhON6Wres
wfEObAi3dwtNHPPBP4xfdobVnLXy8RhG1wcdDsdPJeqJivXK2c27yvRPK0n7sVQc6kc/4CFvd6m3
T5RJ+nfeQA7j9BB7uOZnyUzfF135rBik5paP6A198p7WiV2ZvokGgfEgZdB3bDkCacaDY7h6ycvo
AhRs/FAhfq7VouHBStBGzWenLeTKMdVlGlAilm5ySBA3+OdmrQBX40wCjieJFMXAzYXShBus+K6R
ab24rM62KptIU7RvTqSTlgmNk+ZtLlsi5hq2yHMItoewDZ7JEOMQuEwa/tg2/YX/ASERbzUIUm6z
ffUI7/EE0SwuGouZm+K7iSxjhGPGtGfpcte6WSJem1ZdSiLknP66kHZrMAzS4TPOIgAb6VkPvpAK
vYOcDNDG/1v8d7qkFLvD7/Ek0yI0RhynF4QHMHMriPo+ifU0uEx9lHchxEECFJ2BTAkChF/+oGlT
Cuw/6KCtvv8/3ehCpKPhxVsP8R/qqYVxZ2iFagMBq9NDb3Oh3Glxuk8GiKLbGHgNFHzB04RqURgD
8tzQOwrQkcFq/z1djc9DrcM1cce9A2keP8E3vRmz/ohqA761HSTDSyfJMELo69EBojGoKqEljPX3
Ax6mkDW6WjN6YoI1vhXO+YZ26i2JArM4zd874IJW3wjYvMOhVoQvRRhSv1oP/tX8xIz3gezeR5pD
Lnj0oAtU4OMdvvEYaq1cIJWkfpYGULCqZ0agW0DFSoRYgl0v1J6ije9iOjA8ThvVNRgPC2VHDDVA
UC4Y3tsHiciP6yUaQ4CxxA3ip1Fe2kiGXf2YkHxV/OTL3PvbYiv6nZ/gyDRGKw5MzFgDoRnVTFIp
pCJziwqThL9Vb/5MkzKGtFzkqX6CZvP5aMtMWvMElo6WP58/bUWVRk2P0eYK4Lh1U6mMJ5A35yz7
MgFFn77YyJDPt32Z5jpR2PE5O4mB8nIZ4NRToeWmV1lljHfrqfyYZBAQKmul0GjwSxoPhWirLrx4
XLZUfahNl49CFLSkahcNdKQGtZTg7BN8bOXtRJdcKNcuCZUo912ZnSoTaXF8FowXxyeGghKdbGOW
3vWLz7gJTFDcayqU5qiUeyLdyFsqXOXh34BucAyeCLUa0kYS5CGa/9LE5heLgxblcBPg4S4lp892
zFVo/n4q6a/fctse/oJS3qCvdq92UHR7rk3I+e+xMfIt2toGfg+K0ZAZz/BQUaxNfUDdg0RFAgr9
G0KtXy2p1K20Ck2kZ4XzhOVRu6AEjoDNdTysOsU1NEm5mrBA8s1bIO66aaB4ggnyFYIFIH6XCNAu
yq32KVsCsonIr70hnaZ2rfGSljUWrwLHWXZ+EF56evPNhFFbJ1dby/WIAm3ymX0PLrCjhxpMUrNh
ENrJtbWOPNlNwJ8e+6uOWGv4I2yDQoiVPbYmIty/VX5SKaoOWleCBthvn2iqqUKqbl/92Pykb6ZX
DGpPkmgL+Kw/g55TdXZMv0phDmjiu7is+dKDsasJJLZkQy72W83mxW60FSrD8GLXG4tCzcBk3nUg
/kc1bl15T3e+mG1eTlf3/HubIbzWWkntp0br02Xu+OUUUF3zUV/arOXytSnKKM7NbfsldUCW4IXt
ZmU0Rg55nTmJWbLbBOC7dEEUlOeaoiRpQ2Y8niSUzucWp82FyPBzfFv1IQ0ZW6/o85Yzu9g7+3yz
FXjGKx9PY17stXyapnlvY/9uuFmiGNCW8ld7cNY2C3O9lHg1FpZaiuDVK09UCtpbU0T4I/aKwQ9t
ktLTsJV+scBmZ6F71WpMfMfdB+bEk+oMrcS2rN2MpJWkBf3kTNup7Gny4s37cFmDrKjn6VK7K/bx
L75L6XOaYhLZzMrZOuMEIno0IGEfTptnxNQhZGYraWiAoW/d3dDQRgRvzOTkB4OyBZyiUs11iyZq
+BbHUCHZCmLeIHC6pB5sYlZszanFx/HqDKQ4qzw7yEXoQJQqJhJewubnNph8PPLSiuvZk4lMIbi9
jpKUdJFk2tYzW/OcZoGLnOsJXK87GI+vFFmhQQq7A1B93fva9RflOpu1hNh3Cz5Dt01BSVHFYRA7
55ZNmM/FP/3fA5rbfqqMThMsz51lQGlVk9eK7VSEDusBafVKe/iTax/64T4pt5Ij5usF+IPsHQIi
GsN6X90Exxwb8bwH5nDalywrI1rmS0Na6T9p9EB67QGYCtABIF05uejLG1g3s2UWZ5xpKhKqkcV8
nNikjfr9ypZQvcMgKjb458C1BGq4XxZFalDap/TR89/R44lQMIXxOZjnXl87y2jwxoeutbOkmvAT
vAbHKU9C18Dg4/G+BnL2ro6/U3eW9nQWDdVaHGOaUWv9vKs4PimP+qiabRHA57aNuFrigsAUvU/U
ki5Oi5SraKipWXzyAJtHWuE64MC1ruFw36HkU8fzUdMsbbvMsm6Fl47QXu+mWItX2SAmFr6oJS6W
Zzr8twpPtTiR2L4P7jCEN+dj8BUasOXmCuNQoAVeAzZtNsy1FO8uYPJlzMlbLM84LbmAiv9Zhq5f
3eoYOg6V/W46Tg5GkyTQKCB2nftj6qPpoUAFLDOorvXpIzhxiZZPmjiUFRRpHK4hpTiO0C64Iv8D
yCIv8nl/DoPQ02CH4dLjJm4u6W73qmqvyU51TE2RulDQOdKeZ8UJx9sWXskNAV6pJXMQXH3+xZ1g
fKdrc6mpmRnwGi1VUWRZp5XbDApjr5cLNQkYLy4gdGO81vSuoStNQ0DRkDYuE0YjTdEzzQxm/Bip
dEMpKK4yHJhzbGE1fIT4LMPY92PfGaeeS7NcMpoxtwiLiuPc+ERWlM+VFjricoMxb4Y2VhtDc6+G
NZ5hV3Cbrzl1IF0+eqN7noulWpUcj/Y5tcEwWQCMGBzKzmN869UOgiOm3+I7OBh/pN/b7YX6gaxD
pRZf6+uXiIbAxa26NybKSguU5NmlL3rV56euEMYfklyj3fl/rrMfRQmvDmNqIvtpskf5fPSGA+8y
NpViVJv6iGIi2Xedk7E3+9k66G9EBkFWb6E3VzFyCUdleYBQjuVWW9UO/NbauxBJEWH/4oxK0/7J
l8oLBXwwgX4AMMlknU1bh8Ea4/AG0h+FuUzYKEEryf9iyMayrCMK5jQWADVdyRjkHi4ySus3o3+k
/p6PyHej2x+gEOI2begoIHFtR19Y9PyHHyrEEzdP3eOZoPdy7q7PuZw8/ETQIJW8Nk4fG5iPi6J5
bzYWegRZEZjAp2GQwgRH78kFVSsyD4iK3UfcnBueOybARKrvU0AtsVlRhdt7srL9Uns1kJm5hGpq
pIQQy2+fuO+KyI/I3p+sckZ0IfznK3tN4rXCYUq2HOm7XR9AJGCsbAxjBOAiERNuJVewq917FGJR
tMWfTZ5/AkhVTgk4WwOIpXO3iKW5NBGIjYHOr8UMm33l8ouQtruNVnediARYLx6T17aCj3zwQ9Lb
cSwpls8UcWNRmWVSJGnJVgdYUgo00tZtcGx9tLwUMYZq+5Y64HDhzD9itBrKn7vTM+uZodB7MIJT
iOUbBsMHhfu72WjEdJlA7PMRCC641I0Su2T/G8nnyBkAUOpQrkAODn6bUXOaHDao79EQyeonMgo7
OY/LiyRTYoOkS63d67/Cyr8QKLiEUa+vX/GeYqiSKAvC8IYWdFp2QzKaQ0q+rkFT4S/kJYDk368d
ojn0Y+0F21NEDBlWrZhXtXlRXd/2LNLbSYPw56+hx0/r4BsDpXWyEOUqw70ocgtNreieH4B44mp1
benHAdH68qMknXGwN0hAF/lon3/AczMarSbdTdZvbXzo4mn09DnpNwXc4xtSolyPAlLqQCMb9A66
nqUCatKbIbxRgpVgnQFz6aLfxAojkwHa2kMK+VUyNbGDyg+BCp4q+5pawgyar8mplTSa60Cfm7wN
J1efzDeX3Lu4VKmKbDWRL1A3CaoZRERftBR4ctZhjJDRPsWpHQflmOuw+Wy+Hb+TpSMy0EWg110J
55ST1YebTwXwM8mQ92A6V7/nlcRsX+Buuu2Y9GRSGlFfyK4K+Wyw481kNokm2JubrjJtXAnTlC6c
MFdqcLM9T1J1KFD7JSUvxXc7hzDVKQNdcd3DkRIDAbcAl5n+O7ZBQr4Ru/d5nazu0lGNLkxF2k88
kcsqcCMtis4wYLOvOcF2eUSzfb66PSyvhfZE1E56tuNV+wpZRXYrlc2sa46JtZ3bKz94+JVw4FGZ
qcatZ/PQvZk0FHF0jPjXweIa07MudGehZOi3fm+lzQczADWiPvysnRyBQpUf8pGQBt9qB9azJ0oT
rkO374fSvGdqGlsn0T+YDpzUidizNw62FsJZbj6yKEv5H9xoAgNo8uS+US3CSZL3IOECOHdK7mgd
3ZRCo4hvufeY8yVWHKehswdv36G85ty2Z+qF/Lsg+azRqSsPmvEqGbLAAWNtOo0XLE59zclzt2bm
1AjdmdD3X5S1NTHvOlgbOUIc1fUVuKgDbxjH789mJShuYDHFASZFG9Vlp8o96AUzVRndjLeK/tnS
ewBHHxqDRvpEmsaD8r4J5ptI4zqjUI9wZbctbwHx7gK5QA+bCOAxKqy9pPfkkXmnKhWOJMFVqNgX
n5e+rGuE5IRmdkH7piO1w+EOWKS1XiYS9WbMr8U+zuZFbpB9wSD3vwpy3Zv6rI5KPgZmKPvpHt0f
nvfSlaFQ9zSdDwRIsCl85+YKeWVcUh6L5MFeyTdhdAtzG3gbWVTki9Imlug6UHmztOBKjtAu14vY
myYY2NfFs66+/wdA+tWqX0Oy1TH98+OuW/2o13zYstbRvu0oKdExwhDusftZPgq5eGik93S8bXql
EnzSlk8SN/OcUqNyRUQL3VRNgpKn/ek2k3Mganh9KeMgXg5bMqv2eUn/eE92AhDbXtP242DNRzSZ
ORpRdKNx1DiTpkL6OTdiT6EhuMIWmIu1qlIEWHH4/AGJu2hb1SZ+mi1J5LFF27tjWLx6TpmEkqDK
Cu7sgxXH63+d7KSb9RxoYFOM5ucKJ29N73Psu4a65/DMhjuwKb1fwUCtO0BlB4CmbjsP98mohDP0
76VNtaTs6KvL9pMRIRAPLtpHS5L6f6tFiL3U+ZQF1hKPTDrHmVBVJPdCf+u00lMAPwJvHJ6sAtaI
oVYtl4FGTzzUCXXRWDJHsThUM0jkcjUzHv4UzmdWDC+UY2Dj+Ti+YKlFqB0iy4puYlWAl6ZhYces
K+iBE+DCqB5xRnvHBobSWoa7dXss2gcJNJKKjay8K40RvsxCquz1CQ+OCqWv8IhjpGZItNbZEJ/o
ST/p95JEajJwtLb0XdIGZDUlhBVSYUkZNwt7ecZWPhP7WADBm+9ZXwyX6nV6I75/dbPYvFRX3H5j
PFoqkkkjXOWk31VET/BZkos9heVod3twdM76qGvY4kUOBRHn6/z0UbpPu6VyWZBy+npNAWV5pkvo
e+CgF6I50uEJC2rPcH4+sSdN7rXXLDlDxpsCC9LrorD23d7N9mFS9Avx/zpDLGroc+JkMWAOCa5Y
IdB1TkqzqknmcsRVBKHgGuyJDJDKEpvSXqokTYdAyJFiwL5cJcxDIsKIRvSzrcsTCNr3Cdc5g+C4
cxnNnWmG6YLB94LwEgzBFIMH83soweulbV4kGOHNV2lv/bjE5Id51inuqSjb41LGBOoMiQEDjGrO
FEtvFtjlWWgzSlbaYEgymp3QeY0TroaAN+MhqEScVIcK4GEdcEpEkyaFx9K6sCqFCHkBcOQHtbPz
m+t/rRJnfQrtfPmi5JgKgGSccGHq/K8JL/txTr2EybnsToahpfacdIzCqsNnzehcb1p2/KVOu3VA
4Cdw59DtXKihg/81edXvcxPBoQdeLZ8cd/kAUTcGQZ7vBqFmBNCq5weEIquDZ2pySE79GWAJ31Us
x77wYXK5Igc2hNkQOabtOROYAWzRgbKxLR9SQyD0bZrwup1CEKVXkgGBaGdOs51Ru/3hP7RgvXQ9
QFSh4ZByTej1+RrdXrW++Yt+9vh4EFJZkFlyluh2QRFU9kSRQyONs3zwuBYxe3wS2E6+ZUpuZRaX
ny/JhjY2XNbkuWpt8KySKNBV8iyCdmiqHZZy5ckS1IAM0yCJraXgjH6jJ0nLQuykWoeT0POHub7c
xvSMh3J+rLQ2+2x8T0h+DF3qwkR41BB1ulzT1trGsbGTmId/uKkL3oMOiQqf2X0ExxJQUaub3aEV
SWJk1R1Nw19l8DQ+5KWIFhiM/eZOlnefKruSDS6qKN4X1HaJ8BYHegMpOAQPCDOKOAThX4o2VtLb
ku3pQg1jSyvQeTwoVXVYRTSbaPYysxTY70iBZ/XT1ajAXt14CmjByy2IXwe3g6hWUA6csZkZNQ0L
5h/Fl7D7Z7F0mitZFqFck2ThrjWi7cMpc8NFmFyNM6uGvmJkCNxHJjmKDN+bdX118q7YyE2llP/P
ADC3GhgHOCaGIqMCtZY0KmM8G7NXtmHs7sjYqTeV6d4JgA4ZbJXE6pX3sXSI3NsXceW9a169jnz1
k4Wlx3nUDnFOQ86zDeD0yVPHa2s7EBWPTG+7CLxrHufh5FyaDJX7akadvHDSrccaL0nuo+yfidRC
yy7lGorKImYnRyIlY5ezBr5fBjofRla76JfCnwI/imoDKtm1M3WzT2QkfD88ZRYqNWmqiZLqUd2t
saQHRNc6ZkFAlxqp/kkAjymebCqPa5NZCv+Z96/sOpaT81IW3q8lBIRl+niOA9rquQFghjVc7rrG
LYFU6P3STp2n9P9SGjM2+4W+NzRfbRPhA6NmoPo9PIgKG2DsudIJSwblhxxlhauOGPgNeydFU/xc
u8SW/FrPTCxCB/FLcJqjE3rpJfQM97KvR0CYnV71UjZogjg16ZCtXBEltDNe1hoEpgFNxb0ur/PB
SA6grs79j1ntePozurHBGg+j7z4eP2RYNXl8Sp9VbLuEhv9oOASstvoaf8lDBK9VhUkRh8zshp9h
D2Sya0MrHb9HImY2VXu8D7GGk8RsRrq1/PNofNy6sJTDXbQekUux0Qo7aq8yf9nkOdQ6mQdnh7s5
e2lCSA7w85InTcTE3x1gkXTZBqFWOoezvWgpVZ/UA4MxVIhxAhkyITatc69MU2kJarMDMPg70UiL
goaRFd3a/aV8HJVb2+bgyB8OJKWkXlXh8GXNf/GUl/3d+8Ov6L7a60kkqeOXhXZFweM0VJvIwfO8
ECwna4gf9lydBNgzU7LEtyURaEwQUJaFAj0aAZRtHNtN1IrWJNzLmQ/5jWBrpfCakNJ4F7m5qCJh
C6L8zFVGAOBqaqHoLMz7RM0JJeohNBSCk4A+M8RSfANu4Rz24HcWu92uEWKkkhU6NuT0KSkXN7iH
dAzGkfdiSrnnzo/tWS8M7v/kptvOYNxFwrufLwyDdOfSrjS78uz2F46J04/vejahjxHCjjk8fifx
5NIp/admXLqHBNco3+4iSGtzzkg+xkO2QwPYIrrCXUfN3+lxyYKW4jl8AyOUv0RlxRIqRD26vurz
xa/kEAwz4xk61pt9Inw+pUNY7CZN3H3qK7f13WUYZwm2ffApFJfu1R9a2DTbojl5ax7OKQ5Id3Cl
084AhJ7rEpRLuuDqnkjzVjO4jwmjka7YGO27aXIkvx4K7988SkAFr7bSDrUWMXLGam9yLrdbjYYs
QC1gG1E3/7wmoMgQYp8NvhDz0H2K16mw/CdqzFC024DIBUbzKxtUgPfxCiKDmKyJIWbiB4gZoij4
8C7/Ojc+qFqceR7nU6XXWwdUct2wGrbUuHwqU0GDeElU7b6rIn8GYNRCEalopvYfs+BJObDQ5677
UcWTuDc9htfAxD62zkpnFdb8r+uxcU61t3UONOK+lMLCH+f+ltmKJWC0dWaEalED8cxDZwQ76Pb2
ViIHINDyiWiAItUwhAxxif0RlBzRtFRuNCQzReZvGjT+0t5f+P1ldQqpn8I0NNX5OrjEOUXM2FPA
s0iMpoWQqe7n5CGHXi7DRHfVg0rW6ewah1y1FXBkljlhYusGc0OLR7xEHynQiDeNm84YcgwWwTQb
5YXc04PyPPup7hvJUt2jccrR91wIya2jO1i73roMzjiSpC7rIu+t+W2Pu9X/Efk3ar+3wUD89+mh
0L6KjvvggxYEWeOrVQoNMQSroetvJSktL4ab1q8yE7s7gEMK0n2deSJk+U3Hy1mbLhH78fuGhqan
AgFW671EDErjkiOqLnuOlgo7CRMLWqAZiMCfPDrXlXT10L7bxelbSSAEKfNwW2diUOmtFKhVN4Qe
jmB/ez/8DQtdFul35qr4Qih7DqVExFsrayA3q0B9tnFKXQz4KdwL1fJhCfHea/RIBmptIrnauATM
WyscQJ1+fqQqcCo7k0Lp2vo1xP5MWTN2Bbmea+PMAWVuvR4MlNjlbc4gP6kBv4WBaXj+OWZ615Mo
L22JE6hWO0RjWTZa9dUCfCr/aL2LHZWzeHghfEWQxRaudkdrFtDThY0E2OQUiz001Zqk+hG5UHZF
kyn0HPrjjDefytILO2ixRnKEBFhqQXWDh8Lycj5OlxV+pDUvUgC7EK+wjw4vvDapPC9yL99dWuNl
vzTjpZsw7j3oNQUYIltnfw27XgYRoNgbTmdSVUbu66SXIylqz6KzES4Uir7yO/QWDzZsWs842Mxo
XN96/YSyYlprGcYUvQByagL3tECr8pYdgWT0pXQ20mzba54wLQnsyvBIQNNMiQfsFYCCBSC+QMiP
CodvauNduIWtT+vNSnVR43S9onAeoIXBfwU+TpR1V+k2B486MgtWWO7MgcRImWct6Wy6Dpy3KJsc
1WiLTblQllV0K+3c9SXd5F9NY/ChIaXaHF3uU7z+eYrsjrnNC408xd8jBWBLSgMIgpah3TNJkEdt
g7UgaUGpBCMPvve78cKtf/eHVDmntG40t/Z+VFEFIfba/0gV5Z+0qZfStu8ccnQf2wiGzoJaFsmy
sDEg+K3wCkstSz5RcfuNezl0vEFGMbKJHHRn2PrsWof68ZUuE6QQhpdIzNxXUXfgIuu+F4qYRXhq
zExtd9FnB02zX54hRT/aKgwG8fDtnFMf7XqUshRQ2C/Bpww7Su3wuMtxdepk2heFLSlwvfWusktT
0GCpaDagRCKXxSXa3PJBvtu6ufyd/47/kjqOnC7SMcKuSmCNbrWKSDcaPPVHkxZCAYJB8Q3F6AIF
TWSTpv0a8tynxrcvlhgWgvc+9BxxpFwNkF3l2qRRjiw/1tmV7D12AEQMdYQRJE0MWfpWesNt0HLb
/i99v1jmJlDgs7h1bYD8oy2ADfMkUKlmd+iVff1MAK/C123kJ3bQ8AraEOLwl+48g4wT7VcBADf2
HkeWikJjsBfMIoDJwSjUnQP2MKPK0E39XsmPWI6kcj9amlGxqXBYxmpI/mQ1FoihU6fNe9VWB4Vb
HFfhP9uuFzEnNyLcyFo4xdWQ+kN585g5nQmTDha+nhdczA9sMMp11MfgPAwDY1Zw94xGbR+QagBj
mSWrx+03rRxDyCoecjgMT/4MfRtPB4Doz9mFJIrotzrps+Cuz+aRaMwKJkj2lLIhH4rmJS/wcWW9
LQCNI6kde3x9fuF5iK3cX+8WubVUDDIh8sq/BUDwdUqgzk07gFAmcMaa4UzLbn/Vz0PMVRFiQphF
efvSZs9+NNgIgFYUg/CNA4XQc9Gisea4nKJcZQUOB8StxSF0H8kuCwejUQsNKG73J7cZ+uqbTPch
BYvTnHprp/RcXrAXCCu+qzhHyKmDpxtKpkUhaKpfw0EyHcAglaXe1TKF2fWVr6EwOO6DVE2B+VcH
AGa7O1CBNwp5BwrKl9D/2GmMIgJXY453aH02edr/JTHwKGksNrgEGG6pM1Ed90Q7lUrCyolWfN0C
ZrI5MOs9hReu4BG/Tc1RinJuNFG/ojk3S2bFh7vpuwwm6/w35HwBhKH3LOxYJ+pnjbomc4/SbNN4
9KiurkJl+jCyk4BRNQQ58wYF5j7FIRa6SGx7T4PJVFvFW2xwlEeoUa79FkE9rAxQjhCmkFLWCzMS
sZ6uArmDwxvII6y7/bbwWBxgfAMNX72UcG6Pyk+tNtI8+fdC+88KizDGZRYkyTiFHCIlueM8P47F
KkgWqC8bNrJyzenoPoN3lOrMoPezfl/3OBrmFcpLkv+o6o7bNp6HQ3YmsQU7tiXHZ9nKBtidoToJ
VYJPVTzRSu91/98cjHxySDPfLK9LVdsay37lXDhIYPC6QCtOlYPuwkBmHSKc7xsXxZUu9i4MesQl
afJbUCTqFsXIfS76TrhHzTQ3Kwa/YAZulDOxMKwRE5ZME53w2B2eBdnjbakRKZIacoI8SVkGCZWN
vmUsxTrPDcTlANAneeHn9+ISUbUHkHeLumZUL88Hok9ZibGNbopyjw/k5rndGDd/xjUTZwF1GoyE
da/ZmaKTNaCkVV/F2AHWhCMyPvGY133dR/LYwSm0NKYhlHK3L91VPu0OBlqgeWY2EXh7EF5AF9ES
9p5aJ3/Rpc09/CAY1RE/GbOK717ov/mtezREhiaJdAW+EHFSMepJAvmmq5/i+7qcuBeP4x9LH48k
LoDOO3CwvjE7XeOENXrcA3bvs60CCEaVh8HaLtqxNuriyeQMangx7SMHZcnTLt9/TnoKlUJ4kC70
bqQw0Kh8pKH86eXHIKTyEUJMYtKrLBxr2rOsOzNQ5+CmsoK76uZcLnvpoOAZbHQJ5L8uBxExTdt5
CJQHp0iJgrEuxuAf1grmQeJi5qvFJ1M8HFgokX2q9N/+92N5IY2PnbxeWFi7yA9XRK+D3V/+4VAj
WkfJlT5Np1y21+EenoyCyrBSnKMDeFugovcbSWm0G0oa+nibbKtBhrOCuNh52yVmtrRrbLZAt8w4
AlfIdH0F6AKAmCjbLVbbBX7f51teIofMLHCNwrS/am8SmcjapqTK0WgTd1TITxbifxJIUc5e5ZP4
iGW5fYw8A2ppvuatOXLsExsmitM3QNdsxBymU+8yO/EZ5HGeNXI6CzCpywmJUnYMhOJbkrYsFh19
6UsdSD67wyIs3Ar+GLukp/C5I6Z+Qtd3FP67f3ObGAE4uPdlRzVtRqBM+aKJfU59GrsZsZ8zdoLx
i5AcwclN5MK03dq7DDP6mVFPFMXuw/ivCjlqYeXMKEs9S+CcGF7tnhsF2vcYbnuQlTFyBeVCwZMw
y6Ph6FC0+zMA4oOfcxq+RUpmQgXpSDs6jNjB7hDK92JUednK+vxvUpsk5g1xZjrEb4G+fIjlSynE
itSIfBz8np0nzOw142uX0AtBpHKt32RIWzQtD8HpObnq6Pl4L802SO0W5AKbG+4v+J4HBlcLl+rY
s1WRbePPP8VcELXkKspZnW9Y8JzHzc/Q+ZcQLEiCqEMNTpqEcFc6V4qhSUgY08tnvXRKOL/Nxp30
83RZxRR9ob6T6jtTaQQ61vvMX6tSHFvxZHH+orqYqZfQKH46FltzUybGK0DCAU5tWau5ZNUxg6Vg
ps9VyJl0fyCcJ5g5SEJjKhB8AVZL+uMKdWIQVEDvqOKgDmTvFjHch2QZ4jCeeDslUtPKqOR9TUo+
Vs6uqll84eWGMhHw4Xd2a9lBWWUakQ2LFNre5G8sS9zi2z6P7wIvk+6eaF7Vyx/Aon6sDd4PPeGr
ZTXZnCdeSsQQe22duU81PMdAzsCaSqC3ZWyJ55WruQk7eLDe2yi8x2bOVr/wYPcq9RK2rkDn2vZD
ul1AULXTErFjxTWQsOf3gaBWUB2gpiMbebsgSL3W/dy11bv9XXHChHnbIMIlHIV178euffIUZ4Dk
Dakz7ukg9CTaJEBJi+YRgl7G07lbXiry//sU0jLtETjCFu/nPBZGALiTv/0hRA1J+0joTSzvtmK9
daq0QtZiasFXBTDG2zdjkiXiq5NJrREmB3VLy8OhAChf0XU55nDaPbhKdkYMq7QGUFTJ2EmaJqe3
KIoMpGrYCtL4MDal0OLxiH+OrRmKtDrS2X3LtIFQpy7J950eMx0CxJ7GD5x5CMy3MwzBr2iXumFQ
36IcIY/9QEM3KRIvA1QvcpU7KFRvuK7fnmQ93NU9ciZIMrxVpkTl93jyJizX5Xg9Tchv9pHmkTCP
JnO4DbjFGvUeHamzo2nFJUyvEdA71YCLqq53z215NEGW/LSI4TaQ2uBWg8l48DEhZ/JkPA9Bb9id
AhrNMaTzNe3EPNLIiGUormiZlI2QWMi9x5Fy6KYlcHI/scC6+c+CdQ/HXbmqLXB0QIMCHUZcN2mk
p4PFl9djJXUrniftWliBffosPX2ZgWwfz17S+z2RPRC14IXiBMuqCEcIz1ZwqHXCKvkxpS+8l0yo
sMjXm7Pmmh/59//57OIG5h/T9oodfakqG/N0jQpUyJkHreTQg3xMASf7c2sAotFHTjZdeC5ByF9E
eVcymGxVkjPqx2IQjl0ZV7LEKQa7MjSfPqLFsZuXd4bS2Sd25/jr0TuYwT/jIT3Q8EKv5ycuXXB9
nzob3PQD4QeLEz6s7oJL6/JdIo8LC/J9RAxY+KwXlJ7c/b/yVvoRIHCvjqGCQn8E5Butot1HBJF1
kG2g2vs5DT7C20MrqB0M4/nGMJw2QQmjqdT/bI91gtw59PnB3XTwgZMtQYcoTVA8gewscXMdO4FN
1ooJ6D2Y56GsVKs4Q8s76L2+zI5lWLM5SZX610D0fE1+yiPAAqdHs6lk0hh5yY8qrqppmDf94dwC
xNZrEYHf8fk7RrConmnJ8Zyh1+K7M8l0GpQ2IrvWp/DTnHGtGfF6+vrBzImfprDsXHb04Qh9JKAh
mLWVT5y85gUT/NIULXv6BTieFjjbYJq/7xogh0mw6HIL967rNqMwjJ0xPpqd0rDr8/fRehllEAVK
lX9eoJAzH1wzV7awzSkC+0ODYAitIzs+eaqW2yF/ViPqoyX3//wuPOMHQy7I9e1SYx9dBtMBk1GY
CE9IwPCEdgfSnGrOK0NrfyorTVsBeiWn1OIrZEB98tidUVnkfMzywJUCh9Oyt2LuBBLamhwtlvvt
5S9k3k1CW5GGOf+9tss+uQo3/9yvWAfF0ih+gASWi0VjdUV6AEQQ/bRK7zEnq4lP+tpCfLhbIlp4
bSsdW/QeqkfQUg2VEKEhGKY3oGaw/pvQx1WV2EMKQXZnpFAR/kUuS3fF09WDbiBS3oVs9eR1VCuU
hkYwo903yDKIAJ4OCfLKvWTYALA/V/GTsEdxShJe/LPkuvvfIzHSajlrNdegBgIlm5rFoBOOE2GQ
UQyn9Ow/Q4U8fSTyEt5KDivEt4dCvxyfslltTB+J35Bp74kcEwXkNjosPICQ5b8r8u44I322oe/H
iZJY4tJvDvBJaON6AurZSKtWYT/znTNFXw5dFbJI3azo+OYtd++GV+Lsp0g9DXq5jRV8NM+w2Ivq
3OXrVTcH+qjrGQ1NpLNQlCI/8gGavG9YraRRbRQwMnxw0kgaUadyDyDDYd9L7XNmKluaFF+9IEac
mP71Yh40sce1PIUd9ZDFTMYIbNCeoQtpN8EssrVmGKqBzvC20exBm52wBSBi5TbQ+50YVFtzzaIH
nJj/B8IG+W+ddlsWEyQ3L5l+oeoifN9sF65MqSFWcBM9ZT0EtNpLCkQxb1IL9AOAhY7YZusm9WEV
d2Hqry5p1F5dsFcbF9Cha1mLijJJ+rMA11pkj6MUiZsAoUNo7EIRzL+dtWTSrRpeaOz4ksXBxU9G
nLJ4hkenJfzEJxqHkbh343RUWXavfIZeD/knsKTSlemUG2Wh7DrUP6isHhhyI8seWDChCcR469pQ
nJ/R3z+NpwE2bbLmVfKVU4YJS6O52WbN9JWymucJGdwGmuoFw6UmG1NfW4cw4N+iGQaJE8La+x/w
F71EwKyJao131Ymv4Yow46fnedKGzcbhyu4uGUFLBOYNiqTXLVAE6Rqlh3wmgErqlwkxcHpZ2yN2
IyPVM+A90eOvML0oem5Sq6Tz5xpa1xc0vyz3QG3WOA1s3m9pKJP3CGdEECZN1+3zEOotNTdv9qJP
BI8VBMXCpuShTpD7ElMtHQXCuYu+eiA26qPmN2qabJKSOtRvbYDJHkTJEJlcgR8nrGpqbhhdiZy/
mwNMdncxu45eGmCmBC0V4SaDTG7tIzKeGf0VszEu8/+IlaviqdaBAn79+2iGXNXQxX0ntjrjvWXS
/M3mggqF2T/MVbkY/iKmtwLz7CEGY85BmpgSEsWkw5bsWcQN6Q+M/VUc6MAK+1t3fdXPmggKOZYh
B856RZ+5yXaZX+nduV2geHePxG5f8nGPSeSopgPmxyVIbFVzbHldYhl5My7mKvYboAFacZHXDgwg
L1ybJRP3WMEKQp6wkevvUYoe6hBSWKp7htAOg05ZBhYHmwS7LdxMBuQ0zkOEDTqSdbCUkwQOJnvQ
Mi7LcKeXutgRydNPXlYcd5ZxaZuNmK/3e8ooiu78k3abZqhoQ0nPZz+4OqPHcmQFXor9P5r3f36J
V99NZdQH86eLAmOwvDp2xanvPm5bdIy0k7x/yY75kqVkinItlJrMxrZ6Tjffxg6AaoeBUiEaT43D
u4Ubg+G5bbhdaOG0Hf+r9Zfjx0iRRKiXkG6UVTbdKro9rKLW7GGCWynWxbTgMPeO8FeQaavI8Qqk
+SUnZApgh4vp9aFAeC8CMrbWxpvvBLUlvhfzGkB+tgfB6/G7Nrn2SuuLcKoMjojqJd7l5jLbUzLR
Z4Hj115kCjAEqVi1Zv9Af8lV+OhSAqGpvn9jhajUr/flMXBZ9ye4KOX2XhZ6MvhSbRMUJrHEbDux
KqGDLqWHGcNxD4T1fdoSbI7ArFj2L48SISuOKWTHN/ttct5hQr3bIqjF2buR2yV9hU222Zt60/5L
cH0N1G8uCDu4bFZ6b2ZBME8P44D2SkWKS9Kn+TOJAnPwFuwsst5Ig+t0YYRAsDQ2gpdmsgw7Q2X1
gDYIRUdL5wf/SCqg4Nc0KQVb6y59MSY6dCzmzhZmz4DPvZzW5YNYK8KDS3wopQqnAUj/9EmsuR3K
8ILaC2ZJHcJUK/p0BpF8LkNMmlrVQ6svv3igIaEnSUS48x7tL7QreiQLojjHdOTxqgRd2Xo1xmGg
apTuiN/8kqMcS8fFlg0xG9Iwsii4QYqhvNeUWVIXR/EPt8VmOfdyz/5Ed6PGsMsSkIx+V7F+cGrN
zmcV8ga6P953+YYBarX1raZ2ZTN4KEX/+cLIPWPmyEY9pgfXZSLui58aO7UJrZQ/1KVr5TTEb3WA
l/H089EFs02X74hDFbsHarZBoxA1RAub5SBWDuuNQ2+znJLZCNFbNcWEo/Bcq9C4MErlGmAwiD1I
Gf82UK5aXpCJvyAaQkzRat3hx4mS0ewac++Ln+h7j9zE5ut9FvA1bMX1J6aqJE9lIFtsKTQEcnf2
GcQlaKnGGIzt+ylV+t6t1JnD09WIk3YQOTN4aIqIhvB+vbIL1rCobPX+Nuq0VI11/qdwmcsHwFqC
oRYJPucWPcUcedIiGWGY+9bCbEUS5ZUQmp53wD4HbDi/tJUaH5EKxY1fiq6D9q8ElPCe0+Km/vNW
1q4yIAjait4Pbl6IQcjR6N+/BAkzLlmVkbn6Hmw+OR4iHUJYTD1B71OTOF0Mr/BEIxrqu+4kKJuP
BZiZQbqXI1FsoP+Z8Uzeewl8AcvbDf/J6W+MsuXRaM7Cfm/8ERvCakiWyBluTCoez/sc4cQUVZkV
7O6MGJkA4Gsjh5NR9rJXYb/7Jm/un2n8boRjuk9LX4i3dDkkafPYPoZ02oXG9F78gRJ3SqaFzthh
o5pIngXjoC6CTD6yN6DbNVbsmnbbQG/wG4UJwMqLME1VmzVp/dpAzxE5Xp/zzeCO7hH2R1tGpCTZ
WuxokmT7o6xrKyhRqIVl0/bupDOw7H8Yb3Y38pBfr2Wu05gw9HThWcdPUaDoO1Pu1lH/ksR//ogU
+oeMzvsUlMXfcWXsqJyGepWoY46D27ygdgzL/xpqJFiXC+AP8PEIaM9/ZMDghkwvJWFVDDMH/dgE
fVdO57CKw4ccEQe9QNdGe7/2PF1qoOot/KU8KQmMJv7lC9A6qaOXbtMcLeksHIrns99bQ92RtEaC
bHdUKFBDHGRNAcBzArZ6KnqrMP4pIUMtJCFzFsGCi4tn4Yds8JZ6iogmonKk9+xe0FfR4N0ElcrR
ah06uz4JkidPByehduzRhzWx3jesrAqwW0OK4JglZq3ZKAeyB35a7Z2QOkHYOS60F5enMSTUmwvp
mivptDcXENlhCrFIhrJeLLhhDIkQOeRVvk99Vx4VzrHo8cCEAQgI9XGItxCe8aRS/pvB2ymoL8k5
FcH4Qm26uxp5K3Jf8C3N0Wxr2S5u3ZTxXJwtYP8A1b7f17lFcGHgqXs5VemXjCan9MyKuLNRVsfh
V6hqvkUXvmLG7wikvBGyOjt18YaNJunM9xuvwkvdEevKTwH8aTX0pfryz8JLpK2mwvSA7WWRRw32
swy/HM+tJ0DdP3b/vRG1/5NVl3D+IDGo8I28Q71Tw6CiO5aC21Aqu1QNbt95F4aRhNOxJobkBZMW
XF9Wv8EKAeVTeQrT8Jcw6w20bswhWrjK7lN3UvhlvVW9sohchfa+c568AFVO6c05zRtrOAC+Czpe
n3vh0Y9YgPiqKhPO8C+IvcozbYGmwdaZXxyuh/Ubkpp7bZuBrIZ5UcUycDCqDID1i2lXXwg+XF56
YzlHUe1cs55glNFH5kSCp5MVSj+dV5XxhYU2C0KYwaoxXM9zV+LEUdNQaggVHt87ivOVJMpKOhW1
hH80+L9a7Za4pzETjOAd9GqU2QiIuMmtvOYni4auIViyPRKNxMRbGEM6oHHPhuB6oTgl2t4QLS2R
875OmQd1zZwzcjqSwshpuznNx4obi9qEHAnWYtIuxCXcAVuXzBkkTaJ6GuxJ+7gl+AW8AyAWv0ww
+orW3u33PKVdVjerALVJw5+byW/Cp/iRaCMiGN/R9b6jfqexb+jSnrig+L9SVvvclcprgLXp+KuP
txl2yenHOJRq3y9asnajSJ6wZVwA8YYtd6eTVdTLWkfo4ZOEaccze5jbKeY6Jr6LeOU+YtsAZcez
mjHrwhqzca3yu+nLQa0EhPr2BIuOjD8PhxOaQYVVCEOoc2p4Ve9SDCOHxmccqu1MpmJUbudPY09x
/9Q8Pc3eGqP0bfzkdFi6yC6bs+LUWfkdtsXpJCT03H+iTC/X9bcrKlP9vsE7nmSli6B/o0pavtJ9
Q05DTAGHENtnCb1yuziSE0+rKlB8F1Dh52ihlPJ87r5b58oT/4Y/PSKmYbxoBmAHcGyP2fyVMJWA
acHuK4FgnPhAeQml0Gs5X29qGAMJs6+a6/gIFh70xwfqSfNvqfC0IkMPcRz7WcnzJ2wdjCnuA52K
+AXQ/kcgQl58YGAVLLWWAXRMIVyJggTmqqXDFumnypjHrfBmLke0kaL/0ONQnbdIRzgc5L8SO+SG
kRM/eeB3s4icPJbxcJeOTTVyfT1jppp9X1Ws3sIQSkwJBGSEMiAhbWAzQrPQkGE2cq8JW0f16dN6
z6DAIVIiWkPXYVPnUP+2Hg+BLlF8blxLDiVFMjf+OlG4sEl3RRhhfHKVK7/SzFWooFeA8awfpEWY
C6sOMBjMhMsTO7WjTwlHjh8QTcwWX0enorP9lrhwc2mX5ZOAIZuEhyc61tkNbk3nHMpGF1kyffeL
UbpMzkkigT571diZPR/A6hVPvSHEnB9+abZnO+wPFef6Odz2taJ0z5CZg0K7jJ7hO7+IcVANYCbO
VQkPrQebZVIpaWriNjIgdzdCR+EWIhdv9m3WgWi6XUBi7BHgaSelI4/tsym6Imb0zWae6H+tkTw5
XRVMNxa+OaqAwSY3nMsCMhHm+dtEEO+n481AnEunOFkqoWGR00e3HSP0jQw14WpQk/2GRVC5duEB
GeYZURmzPiwPgTg5K1dJE8iPiSD5lywpZzlmi7aTayHppxg0qFJCJTpNkAoRe/fYyF9WwZk8TNnv
FXyHyQRDfrioBfqYbA/9pIBTSP3yhQBWaTxvJ/QjlegLSqWsnc8IMr63g9XGRjrX/Qbtb6KfgsVi
0tIEfPEI2kqLbhZxXieCzasscaq0OlC0SF7Ie5LDHIMkAnxJbxhy8Og3dj8ddR/eby/NG8eNDEuz
JbIxT5nLDbXMwZuMzEuCHnjVDoPDCS7MMgEmw4dMJzyieXJWjBD2hRRV9iUJyivV39IuZx+tRuZh
AFCAECO7SUY/ifCHCDBuRehv+4ddO8qg1DDbA3xGQIcgF5LqZzoHmRkvGRgYc60ONAEVD87jTvXh
t1v6GMqBDNoLthicj75/++pkhc/flmU5lhiq7vIgcMTNJRa2ey6uvUoKhPtK+wKZMMkBi/vhd5E+
ck3J1SkijeYvvBSg+xT2kwKIVHjwHpQYPMdRTDL3QKvXyvxkn46NedzG5tcgq12bt/MC7z6Vu9Ue
zWxJ7+QtdFFl9pU0KCxXHv4OdEqJdlGmgPwfAT7AiNoORkMYXyalqSAI/oUNk/O3K/OrKMWf2fO1
Lk8nQq8CRrVoQbzuC4OJracvRMrvgy/7hWiepPqAk45TQqhX7eL5T22CurzBl2hCfhTTiS57PaaA
zXQMocJy64RaOG2CG9tfUj6i1Fx56IXbNRtded5Q2k+dyIkQbp+ub1Eds4AeiK/70AO/tgTaiUqN
le3K1ifoA2mtnr+B4ZDKlOPHjB0tplBZWj1LdIKNW/L+5oh4gOvUPRFJSzKioQfX959dxIi3iTh7
3hbzvq9PGwee384o2gm2JRh53E/W/WTo49Vs4SE9T9KKVOzxnuyey0ZUFBelN+sSpzh1Ytj/ZTno
w/y/iFw+E6jcvRWLNGVMVCb82y6OJW1r9h1qnylsk3WIfGG2iF5Cs6lMGKoK2yJTfVQn6okDE7Lr
sVcQ8kFHSTvzWtvRto//rMMLD9a7mNAwuVUyubDqFtgMF/BCH4YFneCM0MT0CJBMJKlrazgk4sFK
f6BuRWqpQaEpFL4g3X9iJgE8YHQh3a35e24UwOaE85qRCw2LhVphp1uB0iHIafP6GkTX6GRPqoaZ
vP3fL9PnW+Y+VDq3DL+PZWpWanTF7zwAPZGxBEiuFJqodjUvwO4GPU04gRi/QzyYlc8W6ck3q++5
i2p4b8RHr6+6WI+M7hYyN2k4GGpUcH4MqPafo6rtrLJouosYBjhYqljDZYhpUHBfVTyBJBNqD6vH
lHsavNZiHLhdQxtumTBi8pl7gvEg1en/a2AfdfxdD1FY372aXuwYzWaeB9mhZ7JC57LvOXguSUY0
4fiaoPVnryEJMPDJT2LQJsEKk1hlMXCfu2rjbMnSifp/hWBaIgjWyDyG1paiIjdlOPjlO+5D4Nks
ZX3BTLvEYWSssZqXLU9MGVn4Whur8dULWvEC7z1nKePBjZF0i8Jy6nBi/enrdwLbv+hb+e2lntKe
dtVoPUIyiveQ1wyhsEIHcvq+ZcocQl+Dph+ggADgIxFt+QFVC4kxhzfkbQdgjvumJ99LQ11Bxd9M
FcE8pyclFvwYXPnnq0j28hme7lH07JymNZ1tcUuB4ChCoG1gn1sVYUevvN6UDSkGdRkzzENEQPQi
eliGSpS2UvIroq7nP8ZGh/unD5DWCSLk9dqhQvPDgbN0LFoxhs6KmxewkFiulbRu/ifZaeEBvVIZ
ErN4Ssth0xvVnD1AKnE4ded/VBRX6OJji3bjr2Q2Lt+kIC6+cksTLffqJAy6Ulh+eJ4jez+mE93k
UQgrlW5u88duYnggudpyXRofiPJ/K3Njudb2jbfqYqZmIye2bPZWgqExBSgJFtjHw4eDDcIJ7qG3
RJHbmQzIcXDxf4Dmi+/jACwYO37r9ixeyuR5dVlYeu22RDs4UTf/srHYR0vIqtYJFENI8e9XaGEP
fdscID6HeZRZH2Mn7CA3XmA9lcY+Jh7IpQVG02wTFCeUDncgCcU937oWWbxK6TPqa2ASkHH1iuSD
PrH8xAoZDak2I8BjQizWPQSpAVl0BpVEevyACrNCZCdqPXcdP6i5jAGoQqHhtXr0IdCkvZXXJP7c
6YAWj7o5uNtJkIaXnObYGe6VhrrXnSk9qUeJok3RMIukOSksMSS7T9XlZxJh2MLWO8+iH20tSuqt
MGrLXo73P9mhmMbQ9fKf8zystRBUlpv75DC6ObduxkCFRFB+0krOp7HVqgfHnBayfd2tnrgelPX/
AJMiUrxtK6nKuSsAW57vAPLanQQ1te+PwFqHj4pzs9Pyt+8S1NhvG4eFWl2YdkPWSa25FzHBdM/t
X1rbdpVqnEt8toVHrwiorsAhd4VfqZ7zNqOL2v5nyAXQIAhGfXOXG3Lto1JKZsRRWYYpvrMUxtwN
9bNRaIMgauoUzyGYVXxsa3jNdjjZnFkNGI6ya972nzkrVPBaT0h8/Q8vHklv0/NJryeeSAr+H/yC
VJJAE24590Tw4o7UZ7+9jpn+Dxwl0CKNexfLeSi3x8Ab0hCHnc4FGuFkfVYLwnA8voSm7Y/DwEG+
COWDbQ42uIfapWzt3wKv1VM90T5UlkGhNR2e5Z6nez4xcWs0kFpMqfIsVnMwVRiYRTYxId+Bxuia
M3+EuWcvf8QxqpqI0l1Sa+d68OzzpohPTNzoNZFJzPoHRUZ16xjKoHaKAlD6TLH1tSRAmmiKVfTU
0qSqpjeMFZMYk0Dqi9ZkUfHmfLc5xNZam+CkHx8t/Qpf+Iwylp+UQJFlLbWCQl9TySt5Du2M7ILW
DD7H8gWD5z1ZHjG+52mWAqud60sEu2oI/MXvbfblzd8R7qj2EsuwrPkYVebjl5/UA/rLu31FGPlt
HybTYhAWgliut9kzTUWs5PGz7Q4WVku5uDVg0zEYrFRY/QCdo45kqqmbHXUWU2lBfLbl5KkSuIkf
e/9/Z5IoCJG0qR/YFkD+bHeVpAIt+scHg43iPOrR3vmgpOJTblP5O7n6ROx8TjwtBPEezZNv1jKd
fkzpZLx1aKuPZhSMQU7eTHq6TslfF7nWrdTSzB3kGVkLdENZnhb/g8/oLqTVqgPT23JXO5+WW8b8
HMisKpfkv1D0NqadRG7DTnLTKdal5K/IPGtpfGQXHFU/LdUD08kE9zvnOeawcC/m/YhDEQuiVMGK
1yhxDdtwtJUHdwDuyMoYu1fhFaHlRQ0XQ8jZ3NscMFmrf0LMHIsXefseyygMrnJGAQtFd09Lmk0V
rB2EcOAZF4xYBA/hIjcQADHLGv5JA+Gp4Ngo5I9slPunnikCRAr51oIe8/iQ/rVCiTnW4TAaer9g
APVKW/Y/Mmj3Uoumy1o3l2hbD8h9k6DBI/VDlcQ5L3qMTw/R+ndyrHAqoZ5Ug0l37Xy9camD6y8H
1TstZjxWRxb+UCGgNx1yoELQvTsWJCtGKKIYj+WROZi+dWq7yau7gR+UR1RUq6C11JUPJ99dg0id
SwMEUsejsRxTcsDFQJUhXywnXdUl1vHCcs6MBWPFKk0qbWczAI2wsawHcsFOfzQWXAbsUe2zBGOw
T8OTBzIqAtxy7LxY/P+2Z6G47R7wvmY7RDJaqSKPqtSFVlwgU0C3+wMs3hOJ4/m8MM3LCz01WiVm
d4xiTF9TzExQks9gI2CAz01IeOCYIctPZwz33+2BiLRdbbv+Lq1hvbd81C7bL8nGRqPT2Gv+ROJo
lT8gXQqQLycJpPxIGBmlNfesRdRcZWUdEqM0e8Vm4mBymI2eOasAuo0+HnurR4O4B7eHhWEHQr2/
0Bwz6Pi2zD0SRLAVGQzP0YilIiNncAtfh58XYXAI1D4Ruvz9Rp7AE045kcKyd2Gv9XN2LSGUaORP
EpbH3h8q7m1T0b+syHs37CZ4JyaanUCIbhQE5724F6WHkcpws3LLIEFeR6t0cTaOdOmB+9BxBGtN
w7yG+nj4P6ZU7Nb4LO+6q0pf8xfSWJyKVWeuDPtTDpH/BdKGf4Yd9uO9wvojRWkIZk05Oi0ljEgo
gC8gBXUARv7T5ckQ2wVwK0yPIobdmQAkFe1nZVL1eF+8NkrsW934F1umxuUfiu5cpgierlquX4XD
E5DdF85Sw5AEk1qQ5DOdzxglasLo61A5ePTkfoV2hHXBxd2JTxagmhvunPMmSvKsZOniNTuBWTxn
Nw+RU7mMmAIe27ykWYF5BTP0wEZCZPN+tE9aNO5YMtJVFjzC8apFdiwiw5D6rCVdjDgT9ta9O+6x
DG5loDnk2rixmG7Q1x68bcHY+rjY+E2Ze5ntKeIfHz+78Mct9G+L8A6j3hYCgLMPzllzNz4Wow2X
G27N5BcQby2KpcwfiGN4Jyk987myf4sNaq8hcKL/jfUVPYk2gV/qQCXXicbjatxHWHmh4Ugx8cZs
Ojr60nIehtBBDzz7+XuBQ1qc7iFpKwcswdze67PkKWKvowH8pYVxinaBWw6sfgK8fpGtgJrIdF44
9n05nGU4nSYIqweSBJMfSdoj+tK4dPNrb76QAcJ7Mg0NuOG5nqiPNQ9MFeyFkV29kJUJOXnpC/rX
hp03osaOIlUhBTrDPQxiqXytC/3KJ/rtrbt1fNhosNdAG59Yaa2Y06tdDN53Og5oPIaYyv97Myly
3yGN3IjwFEBf4hhcyrpwe0jno5QIRhSZuLHVpNIxOjGJB7+D2YfXoEBUANbWdwzp6ISm58+rYghh
B8qvT4cE8YaeC5ikU50UcEWk9zCRsbKg6ZIu9E1vLvAlGPJukHPN7QzMrw6U9okp/ZgqiuDfCiaT
sT5gmZIIyaqCJmfRo5R6hn65RIP95900cXN5CKaUG3U0wrvo91tDCGvCKZ37i0j/gv1LeEJP7LBL
e74clFnwba8tjkJ1aHMYDESM+4GGBmU2KKYEOOdfeqddA6fSQMnx0nVBDdoksdiERJU4l27AgNE0
UFvuoGOEAJU9bJakKdHlcyIscrsFOgycpUYIVX7gf4EG9SXOscCi/wyGr9FHlknbvQ7Ontf7T1/1
LgJCoRzSLtv3l2V18rpdRlmP2GzpQaolkxXxfQ20nTFrCQn/Tvt3lnw3eYWde7JapozHzW5p+hOs
amMUMMhl/TZ4TYxI/RtQZQ7qBy71YItVLzvk5690/U2cPbLSPZhm+AAl/4a/feTAnPwJv+fgFj80
S2Qr/buu04pKLbY2KuN7I1i9frX9vyv0liTsJczaf/wxg30pN/dzZCb3zCzqLqbNdnrWOG+fK6wj
RM9hPquy2e0npAtvG3d4V8K2OUjIv/3Cxjpow2pbxD2WAHsioTHCvmeap5bEzX0wsRhD8LiPikkA
iW5TNsoIsATfkzoSrUR7C3kBlCM+Ji17rAkWpOGvGVmTJTvlnVszOscgo/I5UL6LCUhvDedlAvtz
SFxvKnVo7tDOsZvcpfXVoXjyCq64Wce0vqq4syg+KykYYy7ohwuQ4qN4VCWV+xsW4Nd2jGp0PDjr
jcaUzhtMzE8B+fJpav4pz2fSd9VUOOsdStzBKDSCjcci1RTVu12XQicYvxpNYfKaRYeV9x/Dm9wh
1kmeyQqKRUczDkbRnNHgJaAcaxeBGQwrj4mqC1EWCxdw+3ZhCODP+yZ4di1kMv0DXdlSCwvlcFOP
MrSI8D7HOjA35TRlPTx/bv+KweiaiFyZ5FEZQGWOnfEvW47DGef1QOpfMdLoRYeZJvBHh+ONalp0
cMhVCBnmoXvtJ216iuzOVFwHKB1B+efNGQU8Muy+ZctVyi5W4vHq2mQLgnST7y7GvsqHfLlwDAAy
Q2H4Vc9XxvgMImKSDgeiv2RUa0SAK/eRejCUNnmatGOpedxddEgX6MXJ9HqXlffVf4y35R/tKM0s
kJhUQTHh61TT/xDdxYUm9jWidGUQyiZY1HIsVrHInSsE6Z0fi7OJZVIiA4kMrk38FJDuO1dh+dwF
/oWwAlNWap+vrYvtmLG/V3NRh9W1VMr/5z+QrB6kma/JzMd5PYGkakfkjJUYii3BCJp5xCJHei3+
L+OZ9jKjtpAdKRObt2s6TaeCoUkQOVc83oHshEOGK62QdMkpAzETtNj2mPCB15yiedI/bJdMlDHl
5niTCCTRsRsWP3P7Oze1UBiUH9lNnyTJYw+vaoWzs0P4SWp64oLY9Urhd4oH6OAH/suvuwO28iev
lxH39R8ma4YwQudPbxcV0mz77e1MVlWxbAV2EeEv0Dvux6posYLBPYaewlkbnVYcaxHBSGErChlv
0F7k/SfLOBW26gxrVNKP/wq6Dg45iUxiu7PIIoZ5BynA1KC5yI5gKfP1JZmWF+c59PbDHr9Vr93r
QlhmoO8tfwJdg597vxUf3DrVMeYi+z2XRavPUBhZQ6mdbf1FMZ1j3XtKKkg9XmXypYhcTRLP5/Q/
mOZt/wkP6KWXI8KZ3VeJqqDXV3G3t6PLaKozdnKl2/5PQWzFZPYrDYnmcINW0LsiQQfGZjoFCt7N
qAuSotJ2cQaIyr9yHY0JTMypfgyAENpdqcrGCouL9umalMc9PSEiJtsyvKTxkGNcQz3XXYpFdODN
2V+3tX3wXQU/JKhhtkgpj1P+bWyyZANELrLHV9eoo7jWR6O2HDW+CXYk85VbbteUUniPyON2o4lW
TJErHpCLGEWGwzgmcfxvGdAWVWonSfZqHUF/ZL5xrl+kxpmOFaiUTp0Ib9BRib+Le7vWSx5PDFFw
cnRCt4ZF8mEgEZRuPjnc8RjxI54bCJHdqbypwbq96a2vObAxiQEVxFAnSTUZFEfxAyct5ooHdiJ8
x9qVz21K3QvTceFigHLAMdGFSdARanr6wnBoKt7dfHI8P/nzQgqWzfV0LdbnvRn+vkf+LN8pkxMH
S5hJwlo1ysayCS92i1A9LysxCAE76tcr5sjrXBiSy20piOqcD/5cqqam9byf8YgtTS4020YgPkrh
Dr/aOgeqm1YRa3yt0rGvMGZbVXO92Qp12Wc8mZ2usLxtyiA5BS2EHYhzs1V9aopmrqvPWwAn7BCC
sOzT0odMZxRhojlpO8FflN1xHNo7ptCDLP9cTZ3X+H53KWxfrxtijZfVROqz3ZwAOPmXygNlPVVR
XUy7MjGM/4KjueDmFm+W7v4q82bmcD+gzby1kgsG5qqDUIKm8qlCq1gtMtMDyVeGFiGKI69zX1Ry
gZXu0Fu1ZQX1owZY7z7Jgmyd8LoBSLFTU6OPMLw6+Fdg+ll6HuGopTPFK1eoiqDTl0ia0KByz65I
hm0eMQnFx45Eq+E7SBUVNxpeLEDdJw6yZ9CZCr79+MmOtEv6Ukz5gYRkwpmrVaS+/lKVFN8Kzq2T
wLhOm3/a4QMkNlD/gHkO5vdvOX6BV7vQOu9aa70ZBaCtY50Boblc8suZazNncTSbDskXF5/orvP/
myL2sBpnu6Sg8y1FJ2ZfkMVnjFbHDsbObCz/2iEQKEl+qVWC2ivKk23YIdDIc5PLi7KHMV9XCTI0
+0EGTrUpE3i5PhYiiGOjnWvi0htM4rmcESjH3wxCmPoT20R8sM6ZsvzfpYsL8w8XBa/1RioG6i5q
iFmdmfG4lFY5Sjv5E47rG24DWM8pmmLSIcLF1JCwJ0gWoHGE5RU66ncLRl120i16eDaVjX8HHlS7
lr6LUVGBds1/v+peql6rctk2QJjPu9mgakVPF95IGSq1qT7qjR7XkWAxXWqfWBvANAW8jU2ERztX
rUiRvS2DnalLMLJ3PlDKmjsVk1acqV59bxxOp0BwXRuerMgUp5YVnLUP/v0SWbh+cVkIZkDFUCzo
AKuIF/PqJnYoJ72LiXdEzAyvxqbnCB00KCUeU4dk58xSbO61U6C8s1BUsNVmRwlWb96Ua8M/13Cu
cOMleD01oKHuVGoYP5SG4Omd/7IStJH/TuYQ7VJb2NrsU/HU0R8RUWb7qMTOHNxzXHTYgVTnxODf
sxvPrDsGek1zcwqQUu/5YDCzKdn9Q236VO9T8QHrpn2PSBzUj+Zx5NahCJUumRZb5rHGaTiAWZri
wrw5AVKIokP6dKq1QIEwLXsOhkHYqFgS4uOoqHptVqxcfabsck50XuCuARTkRrlyAVnB8h8sK3F/
atjOwpncVg4JNpc51w7N3pVcGyTSCHp147N10K5GBUov4mAZuP4BzFaAauo5cpHymRWz89rForpp
bLeaY+sgqr4+HTQ2+5ujnYdw9+jzkQiSFQnXwWZpYqAwC+xirkRPyI5TZwQTBtDLuAcYKHLbLgqx
IaSfaE/J0wvvNpv9Lt4dCuDUvE6XHI3kuO2OIpDcZqGs5M+/uPJBUrVv5Y4PZgDhZIz0rUudmQT3
BzEo4q/TE2QbIlvr8gZ4OxaWOzLAbjzPGemakUVRg3KW5zOepplfup6qU6IX3k3fWaqRd4ivntnE
iFzmYeTPe7HGAO82fli2dmMyeZicSObL+7fvfk0o1UsavGLlAxOWA3pRwYJLFnEOK3+yCwtMnId+
UfbuddpxLpcTUusU10o7eE4aQQMOaf8WHYFf4Y1q1O3UNaMnTL3YK+RPmUnyjI6RK/5/YNCq8sNH
mXGkvi2ZavCL0znEq7BD4R5y1C4Iqt+UWdBmKk7thQBVo51CkF0Wc+NfJSiEFcPMjRA00H29KHaz
7sUX/YuH2JPD6/l9CapI1jblXbK9CRJCpWLnlKRUvqvMfgdSGtirasbo9jX9P5Y45KHnPVlMYzPg
cfSE1/tn3/jDoqHzQkjR7drtljRoy99eR0LUYjwbejhVjetkAPInJz2r9/TTneIvtzFjm3tVu8DK
DFh1Nodq61PFvLYoR6jQaTRNyJxL/DkSsBCWAW8kTdQni3HnO7+/mzH1t61xtj0hTPhZyntjySUJ
V2ReFZKgj24TkC7wE3gnbNfmX/A/750ZAMHYXaNcaIqPtxdSaCXhH5TBf61Y0/2PRX5XTAens1xm
h+y8FTJ/Sa6CvITgNb9kmq24WT6hxIdS7FK9Zg4F1ZClLQnJ3yoLPDZup2i56QXV8Qcx64li/Ap0
673ZWcQebASWb3pZL7k9Z4LVwKx5jyu0xye2W//fl/0r0xP78Y5diripwaFLnIHw3hg8YNviwCbj
NXoIfQ8TSeL2t++o+/tglwDLWXFWR9jIX2Nj28zeO6zbNg0sZtdPdoDcshuxsCXDxf64SA1lJn+7
PtVnyPUG262Wt2Eb85ZzP3Zyg3dokOr48XIa16e5K1744t0f4VRAoj02AGq1b4qnYW3d93VXrgkR
zxEgqA59Ckz1+FSmQ23QJpik/v6SD8AfuBR1akqFx3LsFilBdMLVujypjAhbae92HlDjJ9baZOpU
WvIE0suP9XweuXaPS35m47rAdI2E+YhvJp11emrqe2aQkjyCvxDjD9nSDFzmBdb2fKRME5Q4lSRI
3G1G68tHW1F6X75MWSO6ioI0/7q9sqgTZwbUAC2mA0RCzb71zbRQz2j6E5QxjcB8oNYMh+OUBmD2
5HzW4CA4U2OshXOInXbz52gh3gQbK5Ass92MpRaoU0tlPUgzPYGclS6rOsbGo6xGvn0qsjnovWyM
Rg7Qt8b2Ae4xd/hjeTfPWnXkhq0A+9NwCD75u/bQaZZd0Bb/8ZkUhjWuwwRN5zHfjB6b2bR/K/hw
SMPxXKRMU+j//Oc1Gpmqtk+yB02MZDNxfqDRZMYewrI1J/svqblgTLNw9uddyWk1NhZ+JbewzzU0
2ltpygmKYpkzSSixPajiLbJkooUttz6bV5AKy/myTXpMDnFpbfGle9K1BwyBGvRRs5A4KzUwiU7w
9+ts7J5TCVF0f7Snetp3cbTSR4JXcCTToAr/Mx3MmvcyCg+v7C8T/rvSJjixtCtmwQlAm5XEaVMU
Vdw0SdFs7XjXDYtrcq1EbNHGdgah6Fat702JwJ69OqdrZRm/kSlcE6BU9fJ+obkL/XQYOgd6/FZa
vdjC3iNnauXuJlO0jylgylOLe1iFj8aAhLlLaN47wSxASxojUj4zAg5rigc9OqdwRFu9eA70LZ1W
ECelCtfgMDGN1UuISAAWE0fPs3YbXVG7HIjcHvQLnxmJEfPKRsLs7wCGXeMyp/its9nInN5j8bn8
nkHLHHnJ8+C4exrXVJzgb8YlE5WEfE89TS5WqxiCsvosmfJdfGr/720u19Xx48Xf3MTI4Sepc+3a
7SPbKSQUL7kdIeB4SGUWRRrKXZyEUZANthzVB4OqIU1nJqKHkmV6Md5QchyUbGlsHFLHXvUZedr1
Gzr5dAZXTQcrXwvRG/RaCEgAz0fSnffX4S1WrWuRjF4ZzVLb7OaXWe73naF0sle1ZwpbZhrQqwEx
tT1El8zJnsGilKJcbL70dRdUMQdTeaHx5HNrMZ0+/oW0amJiWCndDRqjdl1F4RcUpA30nA3ZQ8ob
jE3nnO16SPPWs0/f+YCwY6Icr1UWoRFMXyWHs51tRMkKejPs/S+RK8grGnUzF6oB9UhKvBuIhQLP
BjOJv7rxm2yvGGBvbrK6dW6WtwlVbN1QnvwDR20/Z4aSE6zkpsgP14utFmpSFIAEhVGxPEhOq4WD
nfkx2mofYwL7gE/x9TxHBRv59znuzCvLe/gY6tu1H9OOMBamFJosgpWG84HzyBxnZX0v6Huar2a+
QtVXcRXix9xl+IreTaQkNHCUPLegdj11QO2s87ODy5PJeRqcq5c40v2j+1W3lQnjNv4spWgTCP43
RH2xprmSdDn+UD+99xNfDpiaM+ayoasIPwktWTH6h0F2k9FlrXx5KRw1e/bXwO2qwwdCaY/g6Oew
lQU5EebBCm/d23ikFzqUubCGLCr6XZK32TL10/n6GvVFKAzVyKbOnvi56am1kd7+6PxF6IocPjvV
TUgJjIgKEGvXrzf/3af7qwOzqOizpJ9M+uDv+QWDcH1yWYdoCbMexUwUEmno5b0V4pa+PIsCWQJ3
z2k9AhMgDRaRTXZilDKeD32vLRceM+SCFSRt9S2UGoMKriXhVdR6cS/LEaowZMYWOxkkC9StErSq
Hf0S4NIBRckCbb/yJ2S4wZVCXgRrlIAeyo3DLSZnGq9mngAcB17KbTCud/k2YNxRwwAoKFRHar24
ku6tLurqRiM9lVnZNtiAselT0UeriksaOm7w0Nh0J2G+aFJjURhqrMA0NqMwHuuPxlyXFLGGv6a2
f0tfID3Rk4gLQf4TS2N94Db/zpWxPjH2rZdZBXpuDagotilXCfGjQtEHETwa0Uth/MskQzyX1r5F
STuoi7YUsrt69lFpeG8L8LNTmJfoafU36zxuS0vAkpPk0XP+ddT0xNV9J7xhO8ilospKRR51nVVX
Cc9g4YxazH1o+U0wFvoAeiuB61t/I+ysRo8aicFR6HhtZ1SrhHzL6pf+KuMC9XUfkY8vAiw3mytb
CSta+1dB7RaG394UnaLLm8JKh2q99i5MMbISki9RX6SzAKI2ZXrc5nmV8ldaFRzo2u67gXT79yKn
h/hPgcytui5JRfRYhCcaB3WIIcglDLvsoWj/q9MErc1Jy/RWTkxPkZ5e+PZz823BuGujzwZ1aMWU
LxtgqfQCK7Bzz4V8x9tpVtYnEGb+heJ1LLBPF5XhhXnbltBnoJdhR2TvK66+uSmqqpgl/s9jUTzE
Xs1ujQsscw32SAhEdAdwkNWLDZNk15tvJy/XtZnCFjU9k8A+9HikNCVevzmKustDqsfciHhx5Dwj
JnhLzBi4Y0aCuIxYAjygxhm1MumJfWKpMvdwl5Ex4NNqYhAXKqzM3Iq9hK/ekoy6eoaRLCVbekh5
aVp5ZzTbfcVYJiHiIi8lFwQS6jBzQYue7VJtMp+mr9QD16WXJZVC5oZmQdtiYSricytc1fG0Ei/H
IaLkXADzTmTXjCAXhli5mcdhhwGJbXSwrmdCgIgE/ZIIVDOKdVYgSIue+LFUAHTWRq1MD4VT8pUE
69ZaXdhniWtsnhmX6EVpLRV+0l35tuK09Ty5MK8RvI4uBrWDoobFwOS80064R3I0lwLnpSrraQtN
GlmnKHKntjrQaYGDaoE2pAP1UeyKfohqgR6DAz6cvTFofmN/PUbxuM39vPX7G6Uh03QJoMKGsYdm
Yw3ApUVGy9/G2Qo+iuIeXGlTQLyNa6voa5EykGZr7tN9JVesnWFApqsP4j+zlsdDMBUaLifku5mh
H+3xhZeIYWMTWAJvbSOws/hEVFBEDiGgB6CWxpUmHw4yxl1iP/pWgo5PV04ochrQVxCrB8mTCRg2
gO2YtOwa7l+9VD9N8EAwIcP2My35zJh4XnHjaX3yJYfbYu8tCR4dTl4aUHlT9m0lAy+vLuho6u/5
eSyEzGSnTTixH1uXJEann13W5nZVRKUBqjIfvh2NiFW25wE1UjU8bJW/BHO7pY0U91GyFIs2p+Zf
ILKF48sbN0LKjOmNWw1jL85+IB3TxDUVDmEJwFJwrlMd474vGYXZcYQRkVkdJBntwRXDF+Wy4kJc
36pp0ycSHJZr2Pclc9Agn7J/j8mRHzx4wBlqZQgPj47YMRlb4E4PXywGctNx+Zd9+C2k5QuYnJ9/
mjRlXgwa2kFBc369elMQ6aOzhSVytiBPQLN6Vhgp4olLqjx+mrO5gwwmkTM+XpwmvsKvHrcov+Yg
LIBT/kOhqWoZZ7LnlI94JTA/nRtK67XIIaBzBooeJ26Jnl6voCcrU3lEwbNOJ/MgFvnY81lTmNIZ
VZBb4Dx1fkiKywYDgRcWavL2wNNJ9ltnzdOBExhDPTUFm9YFREfJZw2KPnLdiwX54fgPWQ9Xupp/
s3a3dtWJelJgsVK7k3rCUHGwbQE9mjZJj8FohyJPkW4LGXOwsxtkTx8BJhvYiGvnXf5LoN/ZBt+t
JvR1O7VWFehXaz5gHxhOvtZcMLvdZfHNVRy3ptkELvttzmGhUnpkOQp569hFAIc1tsrNkpJ6Vmk7
eM1qoKuWsQssPO2s5L4JqzfzHFlwqyW2yBvFEOnfTO05PguQy33RquChmegAVgRHLMI7DHRf30hJ
3CoPQxmyhpcmmM4NZtUhh2yAUDX+7tVnQ+8gjZHes5oknVjZiBQquRtubeJOOAHCiGJOVZ0rvaye
iPE2/6uruBzhs1b/9rBfwR7I+H49WKaoUFjPJvIe6Ar76lCEGhRbO0woxLZOxyqGCbp+MdGjbffZ
PLzOJtc6YugokC3iT3+Sa0mi6LWFp14wGr5TioBG7fKnsz+AwxM580N7GSkmUahHenOg7BN8HXIt
CsaNjrip0MP40lUhbni3NM+mFNTeN02ACsJlTWqTtweq1LDmLSCG7jZrb3QIw/Pu3M8vbOuKuFmN
vRwiExIFJWS1rmxcty392v0jblmg6Ufi5OSrsYO45am2paOWGjgNDvghqCuR5nre1yJPtJBr8yGN
hJ6VAuz3zU5pMBc+uk+hKRWFMXgWxVkJvJDi6IHpWYUMZpY2Fw/JxPlY9SEAMKAbKnglnNAWyovD
0+yZDLZRq/JiCJk+RDoz1YBNuLp0rO1rmexTQVmo77RrrfNIkv6atlUAafxGGy0ROB2kFoUPlnNB
rflULcPHaa/FCUw+twEDDQOKEkt4M/BBbGQB5pmwhSznc8SVfmh/ByxLpzB6kykZiU5UdMsJpcYZ
ZTqGfnIFqkIm8jpnyhiRV1QgCzOCdKJstV3ZI3wRes2Pb2/zkkeAOMVnKlUiAXumwrFm0hGn7JJ7
JXwqhGWhdebNSpDNbqoHUKDcVj8m9+3OiUR3UWeMj2e7NWa7b7HoUPGHDmIut95XHAbBPcbk03UE
9TuT88SZod5UfEdBUZPPXRXmdyjSq8LE/IR0iN77ftoRi71VqX3XW9j5xqp+9W5rTsWWIeyeoNv0
RqHqsrkLd+1excf+Ahq/07YLaLHZ/XKvfCrGXuzUbfv7TF7Zur5vuTiF4cTgbNPEMbXCQf0vYolT
0CZ/BTfth5M3KbrgvJCUM88YwpPzg6ClMs0911h32hCon5wfTrxHeHGDTK0BhhoPh8nr3bp90xtu
mZWzYP9F1Y9y8BEFDKaYvDdKEbcuJ03etzFbZb8VBgjyz1DDTj5X3CyQDDcLW2fQWrOQNH3KOUJN
Ksza5mvxn7UrSqu0XJlfbzXi0W14H0Og8KbYD/rnl+8tK+kb9uTWVs3f0u/d7JIYxx1Vqh9jX8mL
tG2xQ+Jg5WVuIGIbfRfQXClLhHWj0LJCLI2SkC9rInSMDraOi0lSWScHp5sWSm+T52KS+LnunA+p
cl3jwidZYKMw4DA6SwMUUF17oaIkCoNbg2oGn7LFHQkJmMBwrMQ8Udjf0UoFEFc2p4bdC/CMCTQi
Zg/A4eOcBeL2MU4bpWAd33UUSEJtvpyd2y8QDn1v8Ka7z7Bul84Rhx3lnRzDAkp+OlL75oPJEEzU
WM2FovT9OTY1SMGp5uCqhiKKfb1MdwGy7OCV4rB0HBjRagp1j3POfj/n4kG5bQJNzHfyNR2XqSWE
OvRvt2emgqbfGfv9cshFnHBFyEN1QkhH/aR+ILJwOzID4m0sVIXvyiYXnNtPlRBjGmbDEcfQvGzm
XgglsQdjWqY5pESkdu1B7yeCLOeSqEMi9eEEGBKkBW9birHGXoJoDSFfssWZbrGwhgqGiS/gh8p0
o4ifatzc9NujR6mhzeik6hpkEKPlkiIwDyEC0dIwxFpu67HfNImJLrlS0CBwA1TjyO4MSEsza6Hw
RpfBYk2SqMdoNWNjCYP/yV+Zv+EInG43Fv1wFNCqbJElFPvaDPOKcfdWZZJyydZfUQySR1nv5ixw
8jibfTE7PT0hJgSnc9qUjUQMssAVvLqPw2xQT0Qk0zCp2tcHUyIlbvOL0GCvt1OAxKyEH606tRrV
W5nOMxWYP61ruZbTlf6tXGPA5SX6FI2RWBCa/bqBjTFBmU/W0qUNxRhhj7UXUCpe6ZQHgE0Vo/gc
q8w65T7CLiRbg1joImecT+uOGDf0zyTmm6BmlWzSDSrEUjsxip4TrF1ZW13T2FqZTApVFOG+VNT6
jPGKu6pOlSnEYBBH3IeOdqT5/V3tZq+M59YhF9n28Kw87QnLpE/Yyq3SeRMryI6tzoVtmGhgZBaq
dKzmd3UdUU1LaIjUNt9bnLWEVP7GbPJ8OWc/Mc9CHAl5r7NAPQbo6DOcTNP0auu+E62LJWhaCGO8
a6s7RNdVpTqJpawBIa15I66n5hLR4fjYp7EfKHFkGrBKKX0Jer/ytRt/Zhvs79q53+S1mcJYvi5z
MvbpOaWoDuyDjJy8zZI61q5LSaa+18L5hCW5g6yBolx2Ag1SjKkSLLb1BFB05ieUhVYtyelbr46u
eNKAHN/+XIaXC55OdKPLH0/8m60mcFkW+hUusWsbaAH5AcolcpKy4n2vcFPB62+kj09IigLqk0X8
MhfwR2cNa6OKKYWtB+PJFp4kXrgICxDqXJkZ00baJZ9nQcRACWaxLFXjUBX8vXwBmb3aD+jRKJr+
WPpz6fISXP1tXjyP8xapI/05tGq2XC7qgVsFMFt3fWRr5o8KUTnEjoPgcpHKuvrCcJDAjecQj6xF
NouUPRx/am2zHqxXbG1Jwnrg9lpRUdtVr+HXIjAZkr1ivq0RQxE+Pos3YBpgd2eJZj8aA0Hb9D0I
HFmpSiqJytdtIc97bts8zY+iJbRzOM2snrNDcUWozBgvvPevttjmiVOfKPdzus76aqotPZQJ8QB9
USMvFtsyTBy+vLO8/A4y2Z4uARGfJnBrUyXrdnT2S6Tf5HVx8oghWxlh4MOfeSLbTycapeZ16pGX
Ax6DmqJhURr6xMgkBFtb+sdEJEMoYoa/23TduHlIMSKonhVzE+uLX6bq41gPjjT88aS4RNUGLQm3
p2tGa2YxT80W3oC4cg80VakX86oH2+QRX7woRPURonPie/ufGDDy0veKu87kgZHHMo6xhb5bYSKv
Fy6JJ9vvdU4OlIhBY8HSwXzD4stgyvlb4keo412ZQ6maag27Irfm0dGpbS20ZOIRs+d2RyYC9D3g
d9XrJy8l+uqvO9kaAz7QBe8B3YPdlO9MW64fqMQLDbjeTM8G5eiW51q/UhHps1OnwjsK2Rt258hW
zwYh14uoWGo3G5JfNvpTC2N+QP4nm6JNAYvUBtJrvZB5zM7vwOKtsvxupbcVWz6ICMgqT4NMFv2A
RyxsiL4lrGWSv5NgrpxADM3iIaTGGUdtWmoUvn37N6ZaV62TiORBP2aeZDVybwRHe9HppK7lNvo9
KpOnGmf/DTMOkEnoNnI082GM67FTJ0zF3goX9Ngf5HfJsDgW3wwPeswZMiSHAvlFYpNG6XnNYg0l
dRsjLK8lQufF346kev7z6TIwUV2F9wKonqMrGOgzU0qEd2QPjwDxL+7xY7FOdNZkUHe2jWAb6akB
C9Q9xlzHuR+FVYJVKwjv2ha8z6+CvI74WCPCmKcLOZkrYxde77cMBu58G4WqvrbKif2n3dd0SvSW
Fx+TWn7g/REWLCYGMNc1flTNmapOUjv3YFotqxQ6PnP82w/FE8LP2aDiEA5hT0XxyFKWib0o8Sc0
zli8j8+nSkscfb2aWcK4zQ4lXV66XAkdJK5UYfyKzdGeIoETks58k+G2QOUwRV85dtiroHaP6ZJN
8Bg5QUpS64oW0+DYmeqlGhmqgxzSZUUjus0Guu5Pe+oFzOjZAV15XvpmXVJ4S/fwI+lQ8/+rkSQY
D5unSWbd1DJmcp7AFfdbOjjpKS+1Biw/fgSz1c8WvC2/2E4s9IgF9614rBiXEIW/GRmZYk7EJ7p8
B1STNydp2FXxUL9/+a9a4blbeIJU+VsdtsLgjvrxqYM+mfgvfQ0gmyk/jVlDckGIXsuQfKLqu+Wf
YEjngMw5CXliNgeNEsqlpI4qrtR5H71IJv8C/1AVjBNTMB6jJ1z3y7r09K0AuZCxOqhMjp7iN9TJ
yIqsUGLCpCEt+P7z5ATyuPmD4aiLCfrBksKROzevFavnvgpDlR7zN/X5mcP2dSZdLnQrnIPyQl1h
RRMSP72Da4nsQ13iYlTx+Z6q5/TIvNmcu+wzOly1nutM3nM2EAWsr7M73JAm0dOMyymY7N7t7Hm9
z8KHL2loKwR/JJ/nrGTvgAcmxnH1Qy6vWS3xoW/OcIE4ScjIMZ6+/okNYq3Cl4sD7vTe+iMThytS
SWktenzBtOjHMO24Z3jMXncOSnM9VkGmmfKq5pR72w7636jrI5PSwtB2AEQ6VeYDQxC8JwWRkdoP
3JJm65LSffbSss6Au8nSsmITuEzWqSmmb0UPupG3yD0ER119c8iOeWEy0JATvFcJhvSIEffGQ3b/
8zWGHKYadmif90qZuGyqdlWV8vZHxNgzRudz2O8rBh4lgy5vu9iAqYE82Ex+kjkfEZEQHwuyzvho
4Mbu8thWjDZdue9vPib7Rj+/mabNm5nuKcqUtFHgXcZbjcLA3MFgtSZLyQJDd6sS7gLVD7c+XsTS
F1o7Jn6FmWqXitrvxXR323xQcs8DyIgwRQ3+cca8/cYjvrPoZF2lHnJPmn6cnVCOtP5yf0u7fDtU
+0kJcWkNQrMKKqLurkyVRsPbEoqelsyAu2MAmCvlQsZ1w+EDQFHvwwIQ1waIKqCyZqCVt6oSjWId
UaDh0qeyIZ97Dg33TC9pp5IfsiKUIssq1qBpoii+0SnH+wnD91ex0p1TCq7KpYlK6wLfCQQGF7s3
2M4x6SewxPbPEz0yMMUc16dOGJhRGg26HMiBr89+aslkv86UjStG7mmRVN75ZLeeqDCPkVYF2efe
wDCP6hGJw39piM2dE9Srlh1bBL18H2qQKX3eJVmfp/mGKn0Z4Tw/G8KaOvwxnMXN1YOpZ7JVz8my
Uhfj/JxefOIqrrKqCJoFbjle5uqt5kzV6pDLkxVAqeVVLLj+Gv4gE9R8UeDohwdH2L88aIQ6ZCnT
owGIUTUqKDn9xP1+dFAgdA+oJ552H8XJYrM0VVAYJTgiKKxoukhtn+3Lm/nv1jNrIhYyXenl7fqu
iiaHfvLN8ag3konx9/yBXd09Mbk3g7J9TvH3ylmJ1aOQ2OI0Ib9aU3zKw0OkERvnXBmzMmqWn4UF
VCKE7qMkOE2Kn7oQ1bJXC+j9YXKkC7FTQdshULPxJvvnfElcgtEBhPcJHPkzWwH3Oy54uR8jhH29
r7YbXIzKkRv+eL39hWyXQj/P0EV0zIP3SnMXEePUiSstPBiWN/CQtN9x77drDb+p5VLAaNVPx1v6
CnT9MLF79B9XN+aZlT12mSW5xrvczfGwoMltYQ9XUTWI5jxFhMhCcs+aXxK3/G0Fy2HxIKS7kZzJ
iWRM8ExqidZqiuNUiGsqMMdJFUiGONjz+NUnToIl/IJ8zgEKGM6ex2CO6xhPQCEjGQ5I4SM6ghM/
32/+S6zCb7cB96W1A4+JKkjFqGxNo7vPqZGRp0Ikl7CHSDpr3d+7BVe05nnWysayZvhISb88qmA/
Mvi/6FuAG4HV+kSjok4oI0blN3kvasTIhHtRRyMPVSw1nUqUGyvbxuzisVZHyd2x1FD4iwxHqJgS
8EXoqnXVu2hnBoasU3s5FswSwEuS116BxflQv1qlNwt1GpXJ1QmbI7m0ii71XReRf1lIghLuzWky
1esWyZKJyEtfMVEycyEnJRNTAXaIS0Gcrr8+jmsTIi/kvlu32NrLAYQpQee6wr/badvm7b5O9IL+
XF5YX1W4M+8ZZQkWAllrr5DsH5QrX+MyAYNaSTNhwxgimsKAHS18/J/5G9AN1Mb3o7uppgbofmaL
fHXQbVNACEdgCYkr5VLQfgSWenhtPP+Hs40aXeF3lGLhcsodrI7/OQxdbxV1xSVZj+yYpAXxGXMW
jOAzg57jdVjVHnImNi7i6gBKLP8Vg28lCVPkkREwJcw+NIF9ATfuPJcsAIzV6cZ14U26PVDX0aZj
/1wmONUOg6jGehRuPBmPO9DHMe89kMR/z0dIYV7Xw3k18sLCagMaQMR+LpLOBzvd1T1ipmrC0P2J
5YdvHMnSk0K+v4OVuhonzCYH0vMX1hsnvqmt9qIhUBeUH6ODhlzvq6q7XiusdAYshsa1+8fC0236
re8W/w2J/WMxtBUYSclJ2rMgOSjMg1G3A4Wf42jBdNGW3JeGlIKU0Nt2M1X0Br7O4Z2cGIdgMRKA
J0KsvRhWgrDrn5UOZoVE9MbJgkO1y/b9z79IEpyZexOChZ5i0Sq1JR79TrYRNIxtbVKdTF4mO/JS
Vo+IMWaQ1pW6WyTg5YlkaxDnJfoY4R6dDwAgMZclZ7Y0DWwo2DD+5h3ifzb5aeokqWg9NnUfCNJJ
jjfpnJiuUeqsEeV8+rBNR8W1DEWfHutNPxHDZulrrqKZuowKBdSeCvhiZ7OlRvH9dsUvI6/z2Jh7
ugycM72obW5K3yuimoEETNNnW5fCbLh+y6T1xxsjhlBYG4Pu0AYQxKVYMyLOC2FBBc4NS0deg+tk
ifrVBc4rfhYQ+t3VmtWOH7fcWxCs9j/6Ce/4wTQpAJ1zobjctTwqEi+yAC2Y87YXEBQdn+vvP2gi
ZXRskI2hcli/JNEWkoUv3YUCs7fnvItfGNxi9VPIVTozju1bG/VeDyUCcDY2AR8weFdJjPxVsxYL
/zHx0GJs5dg2oWoslnof9oiGfZmi+2RZjPNmoyCIXlNJzBO5DX6OToPaBapx0JkfvlpZgqeHx+zH
v6kWJ20Ok+55KvIxoEdMMJ2lkbwloCSoOUFpSOUSGFwtpevkcVo1dvsfcenpVmvtuKwdRY4M0Kvz
jMGP0Q6AhOgmjXWT9I7vBLFYn/S9fl4tCDwcCT8Iz2/wa0rYflszRpvUK3cABFdWx7sIKi1o6bE+
Kuz8Y4MLVdr8Zj2F5kZ14EeteUFUKY4JvGLkVhm2poA9sAyM2DDMiEZhjB1zZZJzWz+Q990k0H0Z
V59H1qw/dVrR32tzPd5RbaSC4Na/niGWEi9aYFMXo4Gxy+J7+KQBWveXia+E20BI02AGl9TGCmC2
2RmcnAsgf8lCChBt214k/Dn6aQebF1PFJoW+K9TJKsPY1g0QwPGde8HvhJmW97dyWphUYLlNrfg5
1v3bMf4DkHCyvhq60zipBkWfjDmoGrTWhQorpCeuNaONL2yfOW7yQqEqrMeZDb4OJrkCZCSRCUJV
UBuMQdVcJL4Q04IVjqWkvskRCtBKbd8LH34Fv4xHahomLZLKXLIDP4ytSKR5FiUjJyw9pWxTIqcf
K0Ga5sRywlsAgewI6UNwpL7u0xd77DKPg8fzgNDhJSmKGqXcNH3oh4pI2sjEa//yPhUHCmKS/YmK
ak0a3JEgRrOnghQX6QeGb3j+ACsMa8E+igWkAEgvidUNoYYFqa0JwjMi18mXpAH10ianwsftjMju
ewzBO681DRbMgrLRviorTfGjRBFydf/9Q23ovGTn7F16e1rgaBPO9GH6PUKgp0hmTOdK2LXWeGGp
Jp0/A6QhOIyzWcc6aFpdxnG/FdIt+dqra2fm+TSSsb7dP5OReVBDZTMpXvqTDLCUhyoL9t6MBsCK
eEuoezfpIvilS6GMdeXFrOYteyKA02kiboe1TWTKxIFzwxa7flENHOxyjlBBRY/jsXfloCyVGDCY
TOeskRlRjtQG/AyckM1SVxcbdVGVcIaPhdUX1y7mJD+lOS+XS2KlyIp80mOhms7dPbBC1nmzRxuv
Sg9+vQHu4VT/711pAx+AJLLqTfCwUeBeiP/sSvfzq+UqgEM6McAjFiZNbuSwXiZ1uUsgsyxpASlI
mQATmZ1OUHM36k6uLshjquWKl7u6I3fmr+s66nHBFQDxS7BQHhTLm3F+Q+7eFxWAF8r77Jq8BugL
PRMzXhUiiT+d4H3QcDKTtkqWC/4w6nqjVYJDGAPkjkWgmcp05Jm5gsip8vASJ+iShTIuLgLKYolM
ebhfxZ0Eit5FVrXfUXNGqEN//XWkcDtHHIkPhvAR3B5U35XpxLwIzg2lqPttrmwgZxX6a3Ol4+nK
bBtE6vRHy5lMNGopdgZosbzPOxJRjfSVImi62snOZ/oz4rjlk6lVZeruQJe4nevVHWtflHqvsAvp
d0lXxLDtUssyIZ8QwoZDp1qIF2CTTXEU7R/vUMDpWkm22s+nVYxNxOwsQ/zaEFth49TjM5JWwagw
GovyitDQ+HXosUcgO7B8ygS0LoB0KNgy6Yko/l8/FMltowRE0MH6BYrB0ZdYBTzpjpU/GzGaRZaD
2jqksRzl8vk/pvk/h+JtV1Kik17vxWc9yREkT9w7JLl5wfQGtGz0a2cahB3zJ5XgfOz0Ypq5LMZL
I6INi3BXNPUI6Le79hJBSrBUuDH+RP1tK0GkL0ijzuoFH1GcjvADcoiQ5AV81qkKUkCLMRcR/WWx
DDZDZ3ZVCeLofWHlNagzLbqPG2pKwn97vltstE4MnB8o/zC2Hvx1AYaqKdpgRJvdegTquHHonQ2L
4Mp8tZK6HUECk0o+Yuq8HV1Fr7FUIgSbcSlVxP9WSllQj2Zg9Z7H97HepLKfnKe2dI8rY24xXbnM
GXmt5jn9Mpn6mM2uT9k36n5GgmDIT8IltTOm7BkcBtMS2Pj+EK+SEg3AtFNaZvheHQTD9xK4bqxl
qC9WexjC/OAjeg2MJ+iskt89LFmtS749OdqBkKrMujSl5J1hq3m8aYO3GkBNLkwXgZOPIeAc/v2C
AaswXdRg10SWzHltbv9z0f3AQCjr4HnXoJL5oJPHge7LMoWaY9YUSaWTBaodS39zoWvMYFYPw/YB
Z3ttLNKfMW8I0Mey0xlFvuqoHQ3xoWhBA4m6a8gx9jHRmC5WKPJBiwR2wEul9dxU11Ry+rJoC4Sv
5f20TqPLexXYnYW/ZSgI+swRlW9gmhLx65ObgH9rLBaUXl3Q5EbEzSfRW9Fayqu70Gz4CgRFibXz
SLkBeGD+dnLcqJi8Or8hKtgE+y3chGZJZ6AISpilM29WpLwbYr2rKV48uFPxsH6P8yCnhBactDCL
0ocMRFhyc1BEvh20ryduDOtpdVAx9C68dyDkIO1hX+WHaaMoH9zu2DxmV/tsuix+9BqtSQNUQe55
xhJP2VOVNbfsZxTkzHaX7Chf9KK2kCOFqAKABOPGPsHg6IzYQSdEYhaR7z/h6/EE9qiHpXwdbl7t
+rYpn2edlMuo0BATAQbkzgVfHNdpgph9d3FSsklIJoCwSqs0ocmuQq511TywmTCRwD1VZGiiEppe
Y/8IKq0xnvT8y/OB7EHNrRmCO4HPhBgx7/aKXvkwXKFM/r8ijxLvLsN7kBulDk5L3DcIo+Ih8c0N
9B4j/bXUzrc6BHybu/OwxOcOKttssjpJJFyL0Lfyyv5BDW7FDBI/Nsf9XbEqgo+HBC+Dxn9vgU5P
r5ks/j9TxzQvY33Z+RpKNgTU8K001pURkee5YhothaHdHi6eUzOAF0PhY/PmN9ZDS7+Bmi93DueO
RBOMHlshINoC7SqNVfVx8qv09Z7DA1JRl9bezXkurtrhgNRiKWMuGjxvlwrcx3HOtXkhgbeBQD5p
x26jAKBy6SEj3Hy/72cy+nT/ej5e0vwSeGWc55KIbaV+5E6V87MKSUDmHUDtscC+WTEFk7MlIaX5
0DJC4jKvednZz4joNl7qAlrXJ0twX1qMPLVswlmK0cWc4sRACRmt4vY56uZMDSCW638EdJxfL6Pz
7OVJ8rahCvzx2CnvJvX+4Gq5l8MJoIZgja+NrYft9LmTcfuJfbx4vQn3kpwXNz9Q1gSisljmH7ys
OPvoEpm9CTOzayI1jHhshlchVVoEQfAOa3doXBPCyhADlve/bqwQB4tx10j0OqJ3+1TPoqJUUTtn
/esxR0YjWaj6OBZNMiVoxm+Fa6uYBpoznReEXe1Fg9GWPs7RzVji1PSyoWxvvKEyO3JPnIP3NP++
jgItiPgS9CIdd9NnXeyT4uaMr3AL235spX+fWh9WtlSTLzudM8UqrN3SRZy2kqXCuwfv1wi2+eui
m3VoDHyT1GlYOdfdBrGnIoMgo1oybLDZvWDoX5L7Jd6KdMMxCzX8UC9Te+iv0pvCZXFJNuZdfHcA
cJTLb1pb8aSkZGNwfTnvwynlmMcRA5CoGyJ8WbQzu3GibUNdTf6WT27DA5tI8wKdUWdo59Hkqcec
+hBahMIU24YYarac1fUmA5PTj7mzkqn7POxnVvDmBkz+e8lH8I+w9079kQuARU13LnODrR7/RHGZ
6CM1T9UGj3fKkyGyAloCKYWEMyvtDNmhk/PunHN0wJ4GKyTBtcW8vtdDd2w4H2NFZAq5FTdpyVCT
z4XSRgxV7wPvN2QES84JWJmm93vpmxUMM1/tLqPU+AT/suJD9NSamEEZzvmFMYV5ElXG8mjuzGkm
f7ldNwgAQ28PVyX+hSW7vq/opErtu01+wcVNMXNP2MCt8hIaRGuX+rri5Myr/GBQvLhxvNHMRl7p
2fw8u8BQ31bZxbF8pmOIDDUQEnwYmlHQlzp8q6RLzdzQIHzpecQO8w1GaowuasXo3C5yjKA8Z2K7
e4Usb1lp1CSapLL/ObE7m5VA2QiK4h0Q/cov8w1yIqJT+Pvw0zK8bW8xLfjkkZLozG+drKwDFtRa
ZnTwwIQaj7E4VFLebLAUyFRN4JDa74j5qgGNPFWO7eNI77gsfHv0gHbq7tmeQPmzwPJ+c3/qQajX
43oMcTFiqMqF9ynDcHx38LqYXwx1oG4J36n1naRY+qrbQ5cbpSELsIGX734FGUlTK8moKxX/QZdp
GDw5RRvB+7pZxxz5bZ1kC2Slev7suK3LQBRHQxSyiobP9BA0ol95dRvr+/7m40079ucMJM1CReeE
tbO90lI3QCBAYPjt9H5Ss40oGdqn+iaJ+pRXVt7Fmv8AhlYJcBnWiHwpEFI1Qeecb+puamQyFX2F
w/QkaDltu/ZDUZHWV136Zxz5Uz7afMPUTM5ZqTJx4RknxZ4gELjC0bQcmJFPYhjFblqFysuTzGFA
2cJj8Vq7usjKifwSUEnL32VZryUmxPJZBCRE8f0pHkkM9aVu+cJB/gX9X7Jj2M1V+T0qlFzaLHkI
pCbsrIPFuW/ROPfL/KR7ZBXpvl+y/uTbBVL2iIM0Wv3vj1JU2YIqO5uIB8A4LmTm86JklEoAaCKH
hb3ugBk+yT1aNMnYSHP+HnfcsMSIruqddpiOju7fkirzd+qiOJO5c7W0ZsccBrKIZ70E8dKGaC7R
71u50NcnauW/5JOL1mnEBEs9e7Om7+WnAQaW1vSNRLfExY+C+IvjAqYrCFRY8uGBIB4CbSTedqCG
zfUiBqpS17fCnMDZ+L3WfBXP+Ycs89uhGEr1Tm1+Q+FQX+2XUuD/jKeELI5uOnP/klYRx/pf2erU
euAUnuzRRqbfkukmsD+hHziadal303cPdyx3ds9Za7Y6tZLaNzXsRLVz1s/eMg5OWfWzPfmsmxdH
h/cFat60RktlpHbjsm8YUrdTULx5KY2eIQFOg2fl73FbjGIPn/ikCagc8vrfLYcP54EtSxTDNpKE
9Hdp7iPMVO8yIPbZO8tKmDXLjyz4fncfW8v66Jate0KvBp/kWKsiROFw4U5Fb7BalOpWewYmS4mE
ZhV/xFnYLFxsIDQKOQsgdrCKsye158faW/MFoV4G5p7IMD7V+uC+D0ERYeZX6/9PK6TnhYg6tV9M
Iggx+ON53avTmO8ELT2A4Oj3itiu6XgRStgTMDA5ktHRBcEgSyZcaSmydoVAbgXMBI+Vig4chsYv
XZXBfb1J658sUK38Ah8ymOcNa5MQOQrNQgtOoXrjwkshI/kn9+4PDZAMAiEnFRCEpCLqYgBK49Jj
9nO1toClvCEAljG1udm87APfB4NG/8Ud9vRxWFraYiBWUHii2T023vqbA60lfztJYH4A23rTO3QE
1mc0MbIYZhy4BbeDjAJtlYlU7a1CwkG85lhRLRT+1LhGPSJsBjDoBGm7uoyZuubDojlHJMTGxaCm
Lu1ZRYKYV0RQFP+8R4MKoXD1zENgSTnlXEaSTbw/iBAn2dVT0wyS5Tk2bSBDQdNdRvnEFI+asxtK
iIokxfZxOhOaECXDIxnT3fSqpQkE2VV/ED4KJ5OpFuy/1/D0C3wDTRP+YtFNvWB9UwGSDdqTen8t
W/hCX7rx7I2JeBSKQS/ljOOLW7RSaGzJsCiBKBwCpWQ+ZP1gWvI2NoXxhETEKSDX/dD0zRFj1ir5
t1dMqRfJwcYCMkmLOJwrwvH0iJg9RP+9Qvrdn6QPteFT2h5awqM5hT9JkD9CLMvHpjKIFzQn+HPQ
YxemTljL5SwAfB4kerSmdgFoDUjZFYX9px/erPN1Z8BCg+QEbOCsaQbKJGV1aLni9i4zXswfvjpo
jrahvT8CKHnvZYXn+gK+9abzc1qdlbcEwKqmZW9OzEeumHD2uo4qsHoMMMbPEa65h1gIi2zLMeRh
9c5qNsIf/Zao+tZ5PAexfyDJdcuwhOCBaRBv8DtVOozpz+TNPqx1QNNa2evVCrZYaC2qqvwgZ/5P
286NcWl+nz3Y32zESM0pxiiVLrjTYkImI5XLMKTVuUiKH8SPUux82MYfF+Ow22gROHu8ItK66zT3
iOMPtZdIOJ2A3WQUxCgHkZl14cxESCe2yzXKaDeE0ScxQQUGZ57y6ubX186andZEp6b1Bjxoymod
9TAW7nQjWgItJOa9J2u2WnGSdm16PqNiaS+8NYerbK4/i9HiMmNH/kAgppQmwfsISUJkIq8g1P5d
YCBtBzg9plKY6mpdt6aNgHuNvCL61cD9oE5JShbqZh/llr1isosCqy4cT3e21hEEZU+8PmmKso9f
NQ/YPlJ908p+L6K2BHf6xFFlrB5o8KzJIVL8/AbTGlN9T+063RGRJTSWbz2s+L7htLL497mZdGl6
L1nLeKbrZh+K4U0VuliDl1MxeCPHTEks5lurFbsqjxWhRkReOU+a1jFfpf5n01j2rwJgzxzXHrOA
7SkhV2I8Cb+Ruv9Q4kQ1TafCc23vhywA9k4WQVbtYeXFw1QExyPsCSxkXqOAxiD3TBrgNwb/vmwg
OOhL6hP5mI2bCCe+r8+xAxPqNOek/HUbpwQ0l/IdUMDKwnmuR5Twc92iZJUCGJp3rE3/Kf7JbjAE
HjrChnbDidnhZ6WeZBwo8Y19JnC+HZjzceZvFjnoeQQeofqdJpV7Q3xV08y7EZQ2Pu3uubKkeO+4
06UFv9qy2DXBC3JEAR6jdYz5UGqEpr/sv6rGqnWhUtiGqGJteDWyelSGm0qBNhD6Bgu+J4EvHFvy
Ss1x3Lyz6H9sTQ9LKvC/g5PopCe1IK7/bT95HuEXZ4NjGhxDFi5CQ1kJdixDdSbXAoETumluv6Kx
nNc6P5GD0blX/0efnURcms+o8Pux+SkfgGL8/T4Ag78CMHfdodtm0rFTLNwyGvC60lPwRlsdeZTL
lww5910Fi5BxxcAPZyklR3mILlBw4kN540/LsPrL+6cy5zys0TUebEmGiGv73Fr20srlzOmKhcmW
DZzkKIH06sOppc7oJVBk+EEeV/aieR09PDirWidaWU5t+C9s/yF3nNRs+AFSGTFu3aEMahDgyUZr
W96RcLWHoq6VL8djc2Qex2vztbbsf4obMJwNhtzt6JXMIyaCrbmoDs9MLlaQ7FVld/c4Ra9zZoyf
80hCBcnNFZrC+fIP+ErwQZxHK9GbmDFAUSCtdnNUsgaDXNhGuz5WmW0xru8kUguZD1ezHOtopdGt
4FW6tbklSm7B5/oB5cEZ9UTlJcWGWtatod6RXsWd/sIdr+AHJ52uoFkxs2KGhoadqnbeCXCTS/WE
O9E7UbMt6GyJF4rBbl46NZHGYL+OfgOwe3Owl9esLtdyg1SidPSk/9sBRNF+tsiUzzG9mKOjXB2O
Tfn1iWZch1N1mbpFfO/+S20xuvnEnw8xuoh5QKScuCQxZa1n0N3MC16eoUzfn5fiWBaO7V18mcqB
cqernZLFTjuBp9h9vj+DbsK1Hl4E3FPc2tSgeV0XlbX6cF/qhAPNbEzwJsnUsEzn41e84jjjADlA
zB3gnnCT9Ax5CKpwUBTeR32am/4xPBXVGcaFnFU0OpxBcXycIf3O6o5KJPjQ0U7tc6o4PqI8+KvL
YJeizKoTQ4ZR153i04FBSc+SyHj1VklForbg+LjP7gBVcHwPC/ROL783uGPr58ioLGOcsmMyHYOi
UD74fBqGAYk0YU6OY07sIeIv4Fs1g/9wIjUyM1MUnIFaigwY3gnu7KyttEx8Ve3HpGk0P78ZJ+OD
q6q2VxHokLZ+wPBMTa1C1/gpvmMcGNrD9HMNimChGRsQGVAAfi86aWnM36OQBV5tmyuIG55e1boh
oc2/s9gnxZqiZ2x+sNEMjzuiuLz/h19tQgFX0WqXFweShjzSDVOazKjydfDLxFOMWkCTsolpbyHx
HjTojHFzRFQyP2YUJ9K8Ich+mKQ3PUrQndlBwJyplpeE2vtR/t89USxYqZTaQo3cK7gjGwnPMV2p
9nr4U+b2j9tsSARKOGbHYARircmvPnH3W88Pdl/cMd+p6dHgywSg34QG1YsvRaRjmMtBVlisxYhq
0qhuBk4mP5cK1Jqop3fdnepzBMAAoI9NcQtT7uNQ1Ap/Wj5t0Y/4FsG4glSMjruN55FJAz67lgYD
OoRElBTXFn51UyaWEg55pdDlDQl6X7YbCFAIUgKYQaBKfWlapmm2e8hG+SHBT5bE7uiS7QtraHWf
UShPUWuTHTcHznCCGlMD3cI9cojREpR3vCNMrSwjUAdeSxVCGRk7aMqIbMFVP4ZAq5relOUtzE2b
tS+gD/zTqZB56p8z1DdFc8Ek5PS6QrHL41dir+91ebSyOrp/MkyorPxO13z14M8WK+0p2o8kDBwA
zJzlgBzFB1p3m5FZz3kRfnND7/m0FTQJoUqVQ6T3TZrLd88TNaW50k1APo0mM99FwpXh0At8RIGl
5s1j/OXZq9EiKQglfRQpgsUFpB75WmEpPYJpg6tat/G+0CkiAXj+Uh1gHAPeTRGPfoO+3OQNbSTP
32R/C9Hy5zVZrndPnEjZBOFvJolPCdKpTmubOkHynsZ2f6Hsbt6/k3B9cGao+B23H6Q+4krtnJ/5
pQaIYErDmQUbCPsx7ED5pZ4OjI9AzxvdxeRUe7J03S5kqocV9XPHw6uZCAU2wyuLC+Ns/BJlJ4tR
FoVs60J6CA3+pSml55U59oQF5V0zi4ugS4e/Stgk7rQR8pNg6vaMkLNYmyAPEUlyvLdqwU24BqkY
1WTV+wTk5h0JkVHBh5eTD9meyuLeduQof3YV4+z4wJkD1Scc7c9F/4rJJuTdIxxqlv/njqTnvzoo
QK4ZH+P+UjJ0Zn4UKmSAiAddQLn5aPiIFAc5n1iiXesp1YD1JJO33o0ryBIa25c+ZiueZXWWCPRU
9ryqW5XTjlirYAlV7vYtAgSVAHVkfS0cmbAsaukqqW6mpQBVIeaU8NUweVyPpHFGwSS2exn6whHS
Cu7KhwZ7jp9pz7xS1VFXQEq5uOTL+Fi0L8h/joZ70YQOGRn1fJGb6ezXUBwQuacJzCJ80InTkHSy
K/Z92twkdzHpTxsKSDHPY0k0+bhdm07hMoYi7baEV8TiSWi+s+AzxEETf1LUeBQZaMOYCQyohhPP
4DjhjjKBqhWntbb+KHV3kvE0I/58lBWvltHXKbYuRkUK8RJ8JlIUwBMWPswKwX6W8RDz0owK0RQK
+LOtcIQZkQnP12Nb6CDS7Ji8PauvnDKpHANpTPYDR8f9iT0OPuhjIrvC7Nt9klfVJboJGSIy3ZVZ
u7Jk6YsMLH6IYpN52+dWjUkPk4lIrA4z5ATs59obeuEchkIhssMToaSPkRJqJ67Vwsx4oFRGuGnd
8cJN3J17U6+wezjbBjwpgRy/03sCBHnIrV1wV35JqnkoZIFkYfKbZLGXFZSnKlBZos3uQ+TJa1S8
DTQjQU1KM1QZlXDPESF7sY/n8RXOljUnLgCv9PSgj7CfJ2U8fkwrnnN4ohp/FFC4ECMmFS33qsqc
a+AbAa+2yyEdNnNfRRwz4J+ySYaCfhU14JeAKNH8YYO8F+sjN3l0I7/fin8O9k86mIZxxEHaS/ra
Ka4v+T4HJa1Eenp4HIuB2IheiWH7FXIMbcPDCYghVPj+XfxezokQFSETSAj4/v68G3X6G6fVitJd
6PrrndmKXowBrCpz7v36+KtMcHGLsvwmrsWovIzgkd8z8z94B0Y2x0gCPu3Q6lN152acebkm51rq
vB8UOVuVb0wBjhXcpOGEhCboY0FGJ4UEmOkaGf+8W+f7aE3kYIQOJNAWKwq0tMwk23lAV68qL+M/
G7KGJUGkamfG+6hRk22JxMWCJt9As852E4R9RKlQlVjj+nMLpQzWrjWCHa9swIagSB/J05V1VX1k
987J+uSkdFxciX5aGG6zxQdM3GgWsdb9npN0HXCkawl4lAYqbj77fjEXgBuJFU33e8nLl2wNE6HJ
61oauDrbB5AB3Egj9KYQQS2fbb3ikn9ItqGjCE1Nvdpba/0HEEhZ0Dkuc5bQxGPSpRIcNAh3i5tC
SPKC6LUoL2iG4Lb0fYSdUcUmvBxu8lTG2VA5TqHd4X+ZivzGx5F4is3Rl4tIFOTzJ+s1lLNqD7gw
Gntf2r8kxXQnb5u9biH/bzvuIgv8BsefOnknt4sNUjDY0Tgxf8i6y9bWXhnIt1urTfCwuEehiCll
vecRuHh4CE4TTFVmHldJABwrR4k95TITivEADyvqWjZmQm5gzkUcPPmf6JiXyh7rgvnmeBNrgNWz
ABxxtVtQ6DqW+aXSTnHGftT41eNgv8KR9kLtcxvnhcMdRqGAWa3jMI4Axo/Qob/TfOS/Sz/GJ/lI
R+zipsMTqOak4X1e9OY6Sc4CSavwWZC2ARo4zjknTKXJRZV/MVjnQ96W3PayhE+Pwx4EY4MKrhmx
QzVktb4Ov+5tQ7xF5J9mlf76s8NqpYC5KXj16t/ZNsTxcKvg/46pch8qUycIn5VovRc4YqNkcMFe
mBNjoq/2mE5oULTBHBnaINNgsiuyUub9tECb1U94krMCh7JuswFcPyPheMJ2wlOKE6fucq57ZWjA
u8ayhQYR6r5qf2J+yWALdpnDC1Mdt2EZswAPrqNs6zsfDY0SDBnRqeI/nxZPiSAntktFqXCTdOZC
Euk1P+WPZJKIHKLsjQqY4+i0qM2wkSMnSsXhozLVbXY5mpLh2pKFmKwJ2mgf9+RRBnDhL8kK1tVq
4bRvfU3Wpwcd3bK7kR7k9klCNmOrG5Zl2mtW2j3wzbu4kRJUsoRF7ZkyQcAl4k3Rew4BDnmRa8/n
LfY05uqAlz43cEACMeXIvhSaxq7RRUbiDvCIOWnEwgqQOs6gLosDm07sQyWwqcottmSsXk12RRrx
Hu7obsZpbEoP+uhSWD/n2T30ECtXEwhIw5YEhbhdU1hromO3IeiDLMO08dBvnD5J86KIqp34mrXD
kNMEzFWc0xe2SwXNWfDcaLOWjT+NMTsexgwo1Qlsj4VVY2W0RVptMXiMzCPC7l4pjpxNYItTu1tk
J9NUhy44Qs0hi9fwZj5cE+rCejBwWv2NfVz+5bVUsF2Ki03Yu+THjSLT7eM/MyO884q2KsaBfy20
yXlLYQdbl4fqnEO233vgDJQhOuRBCSYIZ1PpNYxyyhC806iVFjlF0yRhWJfeEA6XVLerAaFqpmW9
2qD3IDvwtlVv6WfupndnfzSAjHfEr34RGBmEmH51MGHGUbeD4X/O1Yciuny9TZP4GJzUtzE4JI4J
1LEiFyiWMa2NI82KDqNMZYM3suh+ZrnyFvcO2b9AJKsJd6TsJsbaC939F6fkYfdIdwhjp1HbwY4o
bWat3m71Cov51uyBaYdQPeaqU4qSocxwSuZKiswjdxS0r6FjV5cSLko+TMwRsewVSZcma6SaJZQI
eSXia/L5Zt4NVwOqSWJ1FPq0BO3KnkoNPSSxIFATFnT3wvo+U2GwgOs6keCW55zWWnool8CyInk3
pjNjcP5x5IiNBKlT02H5vpRmzIW+AhtjJYAerwBTtLkUbckYY/vN3y5jPVlc1NYG1gFY5KN1FvZe
CHMMRykNu5Ax8qxnLhVdVE9GnytKOlzxubBboNuwBVxU0UVgiFbZ5vk4FjL1ZiMlX2DdM0MYdJU6
HDIMKY5FTiDQb5ug0CU9c7n+wzMg+8DvVp8R24oNdsYwunUx3mpAoNhDsbA1R5LRsdtTvFZddSWv
0aNl5tkN/mzUpHQE848NksRVLSUX/+AcY6ROWu2ZSMEsr7KV3oJpYnq/n4Vw7Ru01Wfwg/jm6tXD
OMTuXNgrmVIJ1DkufnqoNHCnUMyOec+b5AEBYpPT7k0uGKRGhch6nikAOejGd9Zm2MX9xDkB0HpV
WgqApnO28ASN1LgU8gt/MrXR3NYKx1CCN+a2fyBmEme9eFLVvQKmron6HaJeitPqIMLq4Kk8Wh2X
dorMW1WBnRe8YMph+ad/ARG7y4ifm6DUhJq6WS5CnYxUneV0WSOTQRCm5ohOj8REqjqLQa+djrTF
gSNa7a6VwM3ZiWTtiyA0/zfrYcW/bDjUFb6bAaff2K/mS2nlika69343dbAHUkS9BZtXPtkaS716
kZL19XHVgfeYQ1DQqRLpTRykKaBGBZ7zZOVN6L4C86YhDFId7WuXGLq/T8AxOK6Dl5oJkgSdvD5Q
cc8CwzUVQD6HP2Fut1vIQh8ATHsKj8+7RqMf+pDyQY3dCaHpaNIw747WMSYIpBryzNdCnrw94cjq
9fsO8iMYEGkDSI8BrP8/jyg08SNM337HrrH34Nl9KwcvS2wHHaxmvTq9KQBrMmNO40TyobRHrPtV
s987MxOmixAWrFnO7dcFxKbrcY1hxfm5iCCVY6dp3EB+zMvurnURVSsAOv/xS8k2QNg5IqreHcCS
b+TYk7A5Aa3B5tAwz+8Vi6Lql6yijwmELw0+2d4GW34J3RmPgyXxEHbD+w5p9c1Li1cF560xs0we
wYxl1uX1WIGGABdjiTqV26fjgSlzWzpsTbyIGykoq/k2jD0DKiX+WYX+t67IIfHNuiiB22g8rnGn
5hg2FKj7lKaSJxSaORwSp6lsNnSpbdnoidtcxjpjQNhJhSD8ZfUwIVoTfrxbDoFaU35rOmdELsI3
+osnck8wgxFUrFYuXCv3CHAF1rpBEudffl5V65DyK7jzh1sNdKoc1Vtcg0InuSIfTN+rLChSI9C6
0GTf6KBu0YVPM3QNfn2hLV6x7NwmxfZ5lYxYyE5EDDGhkLF3vaM6MJwZ6sKUWftxfGr5VsuvDo/J
Jx1+oTXfVeT9y0SP07IlF450ZjCh/wCUe12lOGQ4nLqttKPIe3jIUAZMzS/hvuGKrwDk84j8Ha4M
LGQMfqf5ej5ujehbvhpNAcITU7iCHPRry07NQfYKBct2gE7mIO/yiJjjKLmhSAG1fNkabFPhWh3S
SE196EyiPdCGv9ceRUtH3tdRwb1hyQcLcDjFRxby2pwaKrrg87wpbvtC++f4GCdZO8xP5o+7hoMP
LujbvA3qe5GFwsKeWWov1m5edbqQtPYNph8/i9GHSX61ABMqFcSeLwncozPeGAXwrKC5VvwxpM/t
CQcZN2UUynP56gKYvCysnlasnrXsDvIpnHCRrQVts+rP3nBFs8F9cTyGVZ/AxS7RhaCc6x6HYl3u
Fj/XvA+fp8D7cyew+o9FuOkyu6riJb1zf5Z525O0Bq9D6RmnZgpGM9NrS3ntsFKD2TPo5dddVe+P
N/DIhmMs63ebVnBIEPHyZ73e63t7DvkiA3wFST+0CTfAIKcrQDZM8fhVHDJ6qsmIQs5/hzTb3Wlf
rZsuTd3Cj21IDtEWuAKijkM0BfbxWtvyp0xSWO5d/RupJvAeJaJ3gdNTF4Ka7AarT0z0906xwfsb
XdSMxJ2xUdM+QpaIOn1Q4ilO4i/Nf+Hp1IaWh6GDCyGV+x8Eygm3Ldz6YBHrt18RJF2gubCmvgTF
MjndWDX3P3ABpZUJXft1uzS4jffNGV1R1Qk52iaUVjreLuyh+idmLLLvj42+vmUXr5/eyZWUz0P+
PnGhxOZBPR4Vn2v0BHy/vFv8EcOP9UFHatH8G2GNSLfR5Zgi3jKibeUNXBruKt0eVuVq7HD5Qla2
V0LnxV3hyvzWNXm1FkLIrwgzMB8W63GRoQ4I5dflU69WmSawrXx4EjG6oHbdCxPe9wnYSh4BF7Df
urrD/sQNKOa/YsHcfH2hth1oxxQUf0BqQ1U3wzJSNjuI0yHv1QoV6TSBfKllN0v9KhgGIWTUKUv8
MkT0ThtM5fSO/LP64PPmmxpLRuNWEx2lqRYXwgZ9+XeP7tGQcZ2/Y9ZEbo0vohqvxr/GabAPSi5j
SyWGskScCJKO0beOeXU1VgQTj6COAFldGnBE+Mi1Gy+IQruRh7xg2kMPI/Su1JtGxvVL32Hkhk0C
kpZ5NbeVlzDplnL6bT+KYNEc4fjsFIGe2PbnajCFCC4F6BiHirdQdGt8zsIsrYHzt2+7WRtwkuxp
iwbcIYQoyDNKera3YKZQKBiWHFctg6SaJBy/z0ZGYjHxEcUhV58Nr66hwKVt7Cmqrrf/FVGQT7we
Y8vBvOeoT/j7ltJe6HpS7qAASmQXjz5wSRkRAoZj7laWjFwCbNHGveFSaRBlufztHcwqoBBh+zho
TaGvN/pJeMUxezfGCX+e7Qc6X6SbEk6sDFoLAWmOAHViY6bgsLMa1VuoDNaTKwvZVpYbuK1nZTqY
t3AG16l1FKHQn26o+4P9eQ6Qfe0j20U5VQ9BiT8D7FsJpsiuaJBqO1LDQsGHicALU9xUf95v77gh
OdG7Zk6kpJPjQUQuThDYNCbklIhK6ceA43U90q/gvJbgtGk7T9y2nP9CxCZ67eSc1O5/2KFcKwnt
EHVCH5Xugai3B3UloFqzONLyO5OXWNzX/c8xQsWYLDq3OFewCuUaYsJA5sQdAFvLbyM8CG8kgReR
RSwpZQxt+3zTqtcZnmbnUS17J9H3zo8k40hfslwwdCLo72OuviZV8BzgSj8XXS3HwyukESxMS4vH
xrWYK70Ht6UlDtvogiS1BU0v+ihQ1S7yIuE82DdrLT0WLDT9RmSkn2gurwO9/AUkxnnvqkgudYgf
xct3CzNS5WJ7U/m2uLxM0hwroM5Ge32OXWRqc3o6jqOWKxTCFZZHAFamumYLccvYl7PXQQxN2jnr
c6TjM9gV8kdtTnnaFhqrligArzv5UdBPwFL5h3muO5ALcKPNdwfKpTKycgnGNGj6Uav2nsOXQNZA
YW/5HCzQ3L1txy7zwJpoTTxd9v/VpqwQX3Q5XR6QBcHbN/sUaHHRv4ui6d4MDq9mpTu/kTOdCsST
pCpX9lW0AOr+e594xhyhRtiSWsV2xM6Kgu9zGQo5kMtcSaun41jY0mNBUXjcUCjqaJxyziSiuZH1
23lwp2cdoDPyXnUx+Zom3FvbyzlJmXL+aUJZw4zIjdoYmgkOsMhcN60twmrtiVLs26uwy7GJCjWc
3LVlcg6upEIp7efoAOAEOA6B5fZbw930hNswKrC0Y6KmBdI+I+2RAUi/wE6ngVwctIS/52jThYKP
PwyIVTqf2AutD1ZUcz+Ofh5a/quNKqB00iSBqFuLDnFR/pA49ZopQ2IJDatj9EURJn1WjvputC/z
U/1ltSRLgGjEvEbjsBsCgxAcsBLVjdAp9XL4ygaguAvDb1au9JiBPev0bQYFrZiTx3Xy3gMR9X4b
aEpZm6gQItfxLncU4zr4grEUYSJw6hV71GGqrT85Y66dmVQKEgMwQSDe/ma07z3YYVeDvKq4vqHM
zF1nmip4dEfUYvBx5uWLcB/+gdoMKvZUIkCxwvajbebsLFp0iy+KMSCex92VSsUxzQmtrf2Wpb6i
kDlBKBk9ja2lezPuibidUD3pq+1EB44SS7Rw0LwvM+L5WSYA3QKdq+KrxvJhBGAVvl0rSaXR3QeS
2wC7IfT1jy/BkhITqX/wuzfnIWkP63PdJ/DT2P/u+GzyyM0VEggd2EFr4foT3SOQ5ITbq615f8jM
6T2zP83s11/VRlWphIfqA0NkTMcx3GSJgU5fRo+4wwlJogHhSi9bTcPr0dW7bBftelAn07zvxR1W
VnTjoRIhd/Ra7wDKPPcpkYxyVvjv2k5Bv+O5gpHwFJzS35lib8YQyQEq4ixFV9xaXp2f9zObA2U7
H9hBPY8FEgwM1VlhtS6WgWNpz6vc3BLYbNL22jP+QyBnx8lErcfg76+5l/x3zm1TkksSz0/G939+
0YHc/Ub+Xk8SjtiNFGz64NgZJOZNrm61LDv7CTdDi3iu1pBhWRrGpLAJPFKdKDFiwEiRpMYPXBWH
Y2B6fs+Uyk4t5pQHqlI1iv4g84OVk7UALcDbtlR5SZF0JjP3ykZmr7vh+zOgyLDClagF7312qpql
gNmpMTl8iF4wAv2GaH+vTf5kdM6rrF6O+kbh1dnlaV2MUvnAcixIh2Cfx3wmDJ0UG3IdjWtOzq9k
i0dLz8TGfiKNs+SOuh9Q+tqhSJVjSTdZ0yP3UyTQYjH0zVABepv29ZBlC881rk1Pci9p3zQZ00bm
EQSN/PTG44wI+RYrzPHz9lsmWrZsAUXgVDlgkxGJMX3wYFE+MhoOIB+kC3ksNnR/oOhakkQdMeZu
Y1ZDAYHV1TLV9r87v4oFxzD71poM8Qbis4hXD3sBhbGLbnSYf29RKhII0L2t7hlm9cFAqwtvxQn9
frxJxZn0QFFPksg04NqlHaEf5GQoYbM+WdP5Z6Mjcxx5LOEcGM15zXqxgjlyCIGOKAQBSQ9mEHlb
DHeoX2sH9xESehcPq+lcYsHk/yzzTdohtt/XxQDGY4quYPdJ5odEsuxe5+qe5tdnmM0LQUm0tuqn
YzpPRed2cLdzmYtJyplLR+DvR0Pqnu1/Wmn9oDiLgYJjTwKwqwgXkGkY8cffvoaEB4rCUqRzJur6
Ixbp1FaKj4VGHy8LRq6zx0GxmTgdQo0/PLkW4bTGqempEkxBPEx6ypa11k2dfE21w99FJP0yBz0X
f/FYvX3zEC5O90g2iOel6HZejMwGgpJLyW6e4OXS4NSoSNz5uOltHA8WeVn6A6fE/3cHntadnurx
j7k9mL1zNnnAulxrrGlC8ohXLvNxF8arLlyVLKLHgzIx0GFuesYU+6lGs7OqOWCjD1QC+6wCYMt7
POF1JzcsuC6kaIzRYPzZ9lg7h5DwPCEYS4Gm8/zBccsl6ACNH+RFRiRgs+K3vpa0COWDtLyPLi9c
RuzxQ5TlWvXr7WDrAbVxMMmjV26Rxt9S26uCnKaiCNzRgVpKm3LYmJ09BY3CPTKWGPgDRD2heLWu
Lr5uEtMipPZi1aT6aKaYGfhNDbqukCAnNVcJSdbxzPstqd+jF1LN4wtdtcvpayCmJ7VKxrStnuRw
mABdio9KHxb3wnDBABd+AKNOMFNXOSg8uARy60BrwKQQNL7d0hfJyR/4beYY83DiuAuZhOkPYb8O
C2X3oueTVjzlO1TdxkW0rf81vRFvitPm/LaMm1Za9N9ursKyPMwiwTpcTjLEYWdUrbMCiKZ3IOHS
5blCjUOyFZnAMwXeP/MFM5vldp96kITFn5M2UEB+bfWI+SkxK2K0mDpQg236bZk+KbTADR8+e3Bq
VwBw72u52zF5TBzt+kbTNnXKQZhK7qtoNAcJyc0cBglA8gQcCa80d59E1YPtK37kBWpiOLEZ1L6l
7mM+U3EqOM+GFB+HI4NelOg7VbM7pZRLDT5utx0k7j11MXTlhVLe2zqTrX/4J4XIkoXsXqV2HlyH
NPHplAvuAR22gPNz6nhZHeP4x4Z6A8EKrr9yLNSRGBwrFQixPQqRYlNptT7e+a/Z0Rfb308fZajw
mNYCYq2lryBPSwcnPYWJ1qaUNCxv6aN086eMzRoxXjXTqllCo1arS76ka+AysCqtwerkNUGTkcK9
8N22A12XaD6C4OROzhPCGclrW3olyL4NKA480SLRefymaBeeC1T0FsxdRua2jx31Dlkd0QK9towR
pp/JzgaSaspx/tiJV90/ogzKxQzHJWEQw3ciASWchVzf4y6gPrdXwkxHNxUZN1ZY/KsEVItuiWlR
JZKesqtfSklZhuM5+gxI2op5XUen/1rtRwaK0S9LAGAZb8snj01aqnvIEigkJD/4PsJ9hr0C4/Re
ENX0dllDXyHB4Ws/1THwai70Fz6RPd8meDwG7aezKH79YEukN6YR4wHRQaW29FVde1dk6aixrjZy
sDvsUnQty6/JJDi8SOXHmWOro4f3HGOsEPwnAzSQYTqXQMG1YRWWW6Dzp6Tt4SyIWkr+/i73T1Yt
CdGIIl9WbtuOMsGTPWc7q3NKiNyjHXYIUZjw3Vr6vR1680sYts6qROGe1Q6+n3C9cWymxp1rrQa/
ied3rOgWDwmjeLy5UQ9HPgS4XZ4b3yJpr8HuBASMtutj0Ek+h1YCXhDKDkplmGK5W9NhpoAO+YTg
2tSDIEdPuRSG4nbxxOlAlKA6eVwGKq5XsCNvJZKguP7GOluix3TbwxUBDhUk1ENP2HKvK8U/c/74
HAd9KjjXkiYGFuElQb/A6/0jlqscirITEnXq420IU6MuwT4lvYFkYtD1Qa9VmGtwunee6hiBdVt8
B1XLl/gHRPefoURUCpki6yOucuGPgyIPx9qd7PPVoG1F5W3CDw2bqCzT21nW/Wmbrmi9XyNMrWIt
cr5GXkgkU63rCAkuuwbekQ4sUNOZkk2+Fr7Gl235OtKSNLumgfqhGJbamTFbaBV8rT6sYgJ/jUYT
q0bE7mSOleE5m4sSxoZ/uZbIAUyXQ/y++ugIYTD3YPU687N8uAN6lYyf6DpnCZfZaWD2WewCf4ef
NcpHngWw6Bovx8c6EOIffRi949Xts0UHN4KciQV8ZcWyUkBEBJVSjYwy+DQnjkfFiuIVUxQDCyCP
e7EkgQBUMUiwi+0Bjmn3Q9V5QWILBO71l7XyQ6sg5bak2/6xe/Ww4choUrQchXZQR8m/t/fES6Hd
7ZuGQTVoRr5yvYf8i1lJuR8LpxlAm3EKGF5GBSeyUmhL0QJJ+Q+kRmOqTefyHqNRzdxmxuO1RHYV
OyqfgBFePmg+TpiodtwX6ASchFFJNn07R3XWhaP6D8QZbOqWTiUbNV6kZli4NN7NkqIqek3o5yaR
Pu18Uqhi6+aogm56VTkE0ennmcbHOowsPb2pCfWBuVigJdQykhsgbdHE0JXckvj23q5rIMacoVJC
kQtziAVVCFod2ANFHCWDDeuy/+JYN9n6EFzCCGBIqrEy1Gfi8ZiekdupQoBmmVyvob+Jzjn/cYo4
mK3XaqNPZFjgVSnH+6xc1g1KkRvsLe8voG6XL2hXFZXYRa4618+gfWXYLGSN+sgklOdvHwO4oieq
y/Hqsm0hdvuIUkLEdhyr5w1u/xAjHCGhlqLDE49voHhP16XBxxTtKCFGmDG/Z9zIfj0xcNIPwIiW
dz9Co47ibEthPQHNQDewHf6zR/0cFlFxLV4cLrpIkr9grGgUT7W7GKYymDb/CPmrS9LokzL8NA9t
loQ1uk02eVRoXEs6xVat10GFynEYvOKMfU7BecMaRv6MHA2cf8afzuf0UOtALe0vlL+a6MFK5QxM
yXToSSVT+EA3ZDsuumEsOzDzOtLLFtEiPz0b8p2+YY3oG2tLkT7Hl/uIWWjVdMaFK00RY3FSZNXM
Yc1f30aQYra0dnsIobACYhaqqJMIV8/oaoo+5yAwMPk5WlgbxRNYjHYIi9tHIhzetNDdoOiYxTtU
f+aQX6u+IoENKwhnY9r3epEsO9FWMSC5nofOXrxQdhOPObkKQxN6j8gAwuyN4iZCmL7KghHjuBuw
zhJ7gvwtTYqT4fPnvcasTsa/9WGShUi7Sk/FutczbKOwyLS+8696eq03RWmPvEzqJTHUUFtWLYZe
yPkCqdCqzxmFko+uJhybv/3XtLHJjoce2jXDnXNxmksC4tctJjL0BbqAwTvnSD4ogmCQ065bdRAV
UB+oTqO6mf97691/JOlDddr1aKjReF4oUXztcdm6duPm+CSQnbFpVlvzGh8O8N+lG7Ep0erGRVaF
e1U/e01s27vnJGA1yaBZpTLLJuw/SW52ZvIRLcNYzZoaW/LI/405oQnLcnTm0fEkLKW1+pIILgA+
ufPFT6Qf1bS6UXuD/SwUz3IWKaYEh/fI4lNlK5oxhRRYmZYc4+/crW8AOmK4U5uvpYXO1d4yjwSs
VlaFNSxv3AUO+3TEgWHY7Ra1k4k5/QF7noCkhV08iAHiTcn1tEgmxB8WwAJbn7MB6Uf1UntgsGyM
8MBg64bri++BlqDph3X+N7xPnEzTeWeVGKsow2d6X3K3Vr5MGyvDW5Lhk3KsA9sAUDBqYCPFSjuO
03X0rWuKElXWDfP0o6W6C5INH3tBtfOdXFqO841jQF1Fj/eD3FHJt3fl9ZWMKs5wn2RqdCETNgW5
JaVhBRWHAMK97mT+ZAuFpw1Iyra8pokVBlngI0a5zhYrWG9XENPocZoI70iN0SzGuZvG2PNTP1k6
Uf/UQFd43LavP67taE75eD8QlFyxYPsuHDGi2/I4NBxn7HB1VENeSEkIkQmZPqgsSK8wZDgv3FLu
BvPvwG11qDKrFyCnbXfQ0NG6HDdRi0CsnA7OIReayyD7xtDca3a4enxKUHNbZeFX3wHcPzQe5HHF
tj1hAv4y9kWCrR7FxCdPCV80Dm1PZfMGpsCakebqfb2ikns/MHm8+j6BQplYNaOqDZBPI1DZqFKR
+gbURSZKJpoCydZrVRHrV1/HwPlT26gdfaD4OQxGfpIHGE5gr3w2rV4dhNBnG3vY5v5OSzz+1yxu
FiJTDXhlPpwuplAOB9p70aOCWkl7nIcXyIzuDrVIYrUp9Lh4wEnrltIz8FsdhHxF8wFbZnWzoIRo
i40vIqb0cx7TIitkFM2sK07ToNbhYJaYmGf8mjG50i7GvuP8E+AzLkGjpWoEA94y8Lb+7Px900H9
ih4mUMXkdfxAsXWVpSKrZd8Qsqke2XoeEJOViQCDwjV+OSbte0380jhjCIUNhP6eFqCHshKYjqBy
PWUXK/87PhVRicehVOHm+LJf1Fwl4jiZw1lvonws551y/+tLDxWuAoIw2/2IRou9qaNZvm55KRPh
jBPegm6IQ2A8HVbAx4/6VsVmlWKwa0esmb5V+ai0+sJ8HRzu6c7yEim0eBmw5CWklInAUpolsC08
kz7chiz6aDMDjE1Jt1cY29L00H3Lv0rygMymmzvnUUKo1fh9qSSINbz4uP6hFn1OxKVWVk4u3d0r
klLXgG66SVLJL1wIIKNzIcKFxw2hfKxpveWtZrPpHquHr08n49iDRIK2IO4oQN9PJVAXFVoxu2y8
rP3qF2dMZ7t/xbNMA4x/LONgxl8MtDQ57Dtkxehwnai5Q6SW4XXBTHgkXstjFa6Y5/6jWNWmyEoV
1PisKLZBcskWIn1T1buZgF5mOzo8n2FxRhRsl+mV2oG5n4n9/X1o78frRoXIqKFqGp8FB7Qjf3YC
IjWRv3nHRiTQ3/kT4+/9kgaVgud1mqgrNkO4jtzavk9h/mc5RTK6o+bl/HiT61098vsE2e4bsm+S
hzewTjGGDUH7tprqtINhYt1WMezELSMBCDgeOXsYVWjBI3iP3AR5+0lfzHXCz6OCAVzgHk0HmxUG
//qylU2SP9w0tq2fOjv+v1+XCwVeJVVTX4fCVbWIBGRxJrV0jUG7YxHGsFRqHPcMQ0Aqm+5WXLtK
uBTsTMPwqsuNOZUpLx4kzPnSGJCd6vF+QHOswXnFJN2ZGpndEKy2oYRc+4D3WXouNoQTNudcxGIz
UZ/kC0guCBbaRQ3njktrfcClYW5fRNUBaw2iMlhayggWASdWZ5uZAW+Zkyk6sZ+sh5VrG2qQByki
K5Xm+j+JZ6mRPDXm+0wuXtPlBWy9Asxekxm/uLaFxpRvWEa/td/QxTb07YK9iei82NjQMhOmHOLo
kyIMMX9AaappQNbxnY5uTE1GgAz5a+lOQqA48lEwJZ+COHuF2KykoTMD4DaMBbhPlCU73Snj7Uoo
jOVfny95rf0Z4prmtG0xrAmkUdJySGYGMTMtpVwmB9ZAlFk369VwWBZ9DnDCNAs62MAGeSO1C9dZ
Mn9dyQXUc7mcIPGLb+jxuicUqoftsretzZIyXk6BpR+nqu3GHhli3Px7uvLp7m0r6IQ7PJdcTJe0
MXb64KrAGenLAU3xMW6kOez5AN38UMwWnM34uE+tjTYaY7TM8XP58f7DTSNplaYhbUfVy+MCG7V3
txgv+13iY9kqM+2/Q6hT/9ccFINSL5abCFgm87dOkm0/nAvwYD/cODMYNlNZIyf8i66EWxGBZqzj
ZmHlG8em3zmc3n3O82s2faPqn8iqsahHCu8nD5LkcMexPExPwj9/kiC8569xckhW4G4WO/2ZYiXx
PZcOH8DMoSKRU60JO/Nm0JdgGG7nRBcz6Q+DSY0DVubnWjgsr41Pp5HeqRfXlJtUroIS/uQbZV/u
qP7Eht3JE0f7+T5BybHoXhXf6UqF3AZp0s4aafVYzU3zT+fjaVmeEUAswxsKngdgYr2K+NhC09+F
h8MedYblOM7TbR7A9TJjHgLs/H+ui4gNMPlj3dLLh+2FsBUv7hlTC4atVgsO+tFAe4zusD879SyK
B0WbTXEJAK15eb7lcGOodYRcCHCVuRJIJeRuyWLNlfH1vONTanjvKTgqcElTArrgjo3Xh0jwWWlB
qvm7SDymTGRlUlARWZ+RFsfRxi1mXIkvrk5DfQDtgvcNK1377Al9nc0bRYirFnnne+4yJjI5EP6F
tmBPsubTd0VN1/fIq3FuVYqg7DCwFwh7DwPx28w3U1d/puaWqvzvRi2R0ViQorGYrGuMdmNXkaYI
QMJi4gjYAGP1G2XRRNtrKAvaveSzgHAw2bGD7B3NYV/TgIYJSkkZ7sb6kuGaRmDzbUjFkCd8eU1Q
/nU7YD6HIo5YwSmo4PxhoRcBAG0qVUR2HKcA4BWAUgTqz0RM5KhkQLGKRTlg+LVi+XvFL3TlN1x9
jZjZ/gS93rLdv/6sMVuttXsWL9DkquqkZwnHxM6XJGE/mlmmwJ5UAmo6c/hOYgMsQx73MzI8JglI
qJNK2i2rqzoFgr7PoibSZUXf+8z/pG372Uul0kyJHSkHxZcrc18bBuc5kbNuzEBgbnk0Q49H8zys
92NPJ6k6AHEnElNZL5TyDoPLBK0O+FtqxK2jMyq5ATvHJB/SagDvXtkuNdaq1vKZHNnYg2tXJONS
8FO9ZhaLy3ag6KltzdyrEloXl8sq6JBBICpAfhgeJw4YS3o1WcaNsu3oGmPWHHBqg+AccjQaRymz
pO1CPhpFa4fCbqGPBxBuaPFw7rE5bw9hL8S/IkR8GkYLJQRYxTkXRpDYm9MdVGMvFrgXubNlQoq9
Ho3VDL9vkaSbm/W9OBGq37PZxusOGNppL9a6b0iiFwgVWpezF+GgAgxfWoERvIosd40+hrjlqnJ2
1JNZDAJ+q/2jy6VxJJLCAN5XyE15JeLE9pKUD5Nk+F+pY5jU3sm3jVPQ+qW8J81muimoapZYv5yr
fjolZZB5qzLFt8efR2HTre/q7SO4Kp85Y+bOZN4Sj3s2AZ2P6br/NY/IhbD7YPmzBK9qBS6IWtIh
WaxuDWDnF2sbJ7S36zU5QunXwbHaac3EswPRMHhIUfaiUckwxrr2BF2msBBXbCJhjydDXnFzFwkZ
elPQpBpHPmpQPqKHxBVKelZh5R+e1QMyETESzZ6hzZIlVC7MNb590/HbcqcruaA/fO2qBe73EGv0
YEHmnMXkgQz1kTEC6paviyBWmqZwxhMTfTOch5O73tGJ1FtUqIztXgVo7itXV+7VlD2Rt/HLRMG9
mwf7JW98E6pTOuWkFe7roqOM0/6Gz4g1NzPQDx2l8EpaGCHbKG/ziwHicGPEoFV7f18zzGvUWCVY
Nt8Wn5GaUjqSdIPO/izgZBMRdKjPrw82ZkzfgkuN66UeXpKfJbIMYl1Evt8m0dEivalhcs6kvHVA
fWx6Nv7KTbO27Bsnii2u3/CwBqrIFpwdXycOJnIbEN3f7TDo9FtKwW4HHf4XvVuR2vPipfUaX/QP
P7igdrWcXa1ti5ciNK0zuJ8HtXTUHewMiLQUi8FefwNig5adeBbRuJ50CzeWI0n/GwTiBFT0XZ+0
DuyFdJ16Tg9A1gA7nZf4vtav+54PgKpVprRx+2PzN5b7GDr2GIX3GaEiCEPXWarnipqJwKGMIbA4
iJes1gSq5bdrAEHUx1BZ59gltigxmJ9HgtB8PFeBnv5FvJ+YuBzFt+kOTkOLXqIrSOOaRBO2AFIh
JgSPa/MFxNIPMNd82cLdUs0oQtL3sBk8RuEDPb//xXBXEu75MnCZUz++X0VK50xkSbZvvovBDuC/
MJaIVGRRTptL1zrZn6//1eD01dl9U1bITMemX1fPr93QtS0faEAkMqPOsRXcg55vw+p56viE4vrm
baAqu621arCy0E9YApHA3/848YsFLtZQhKcsTt3TOzaBGdI14iKAMTeidWk/FSYs8A1XD3FS2Hx6
4xOsDRMF24vG0yP8II2Pl6vV2B7MNOpC34dSWuIS5yUqC59MnZjrnWZqTKJ4nH6YOdvrtqLugjg9
3gt9bIyJeUugqJqh1ddECxWOVZAmunZ+wi3xHdSh11Kg/JVGxu1HWpk7TZFOZ162T57u8V5fB9fn
8HyHEypuYzLh55bPFg0TzlN1bsI1q+cG2JRcTB32kz0M/x0AiNQjeYeVVu9Hots7Z9fn4k+QNRZM
ObeXBnn8jl9U4kXABXZQtRwKjtO0bwxcehhn4PESlRkgcqaeSiIBQGGsy5bBi1ooTlaa5fFXgbER
zzTILS+/4W4hI/UYJFC0WOHwhQAUhGZStmrpyyHaPr8BYcwkDkgEIplizGgnKcVqS4Tvp7ZmOSUF
cN33Ja5gRSSO1//O/2dNC68XOjPNSl//6awMNCu2m+a8EIp/EI6A7Wg2j7Cu8Lc3iOnzsz6zF2aE
Xm+qv87nEWx9S4bhkr4SiL/lrinMcrNb/YIJIfaZcBQq0KpeVvcrZ4vWXUr01ZzI2VSMWk/4S8Tz
P5hwoMoggnJwzrWudXyK+t8WGAScDOWmhjAcN6fCOypDgHJUIYF3KNMOsJ14nz5GtXf8I0ZNhNM6
jD7yYIcsR3Rl3Izp1HB3fLFlCwp+U7Y0tYn9udK/OYv3j3Xh1suFo59HienrpdiN06s/iaaDJNWe
X1Qi/muv4QrYfofpXvIjKQMhPFwXqFSnb/LAgVHf4exyfc7gGpl/wIQDtqlUerr9bqiz66jJVbue
ZbIJSV9mfwMcjUVfW6KTXg2Z2KUxZDxKXZRCW/bKy5fhzsLjemDw63EAyn1Okd4HKXa1cjpiXSjz
rZu8APWtdCRwq5bJHLTAaZ8nEIETu3a7nk0BxqoH2l18N3sSH3EMoayyogh5i2wEwZAl40XnpPNx
+l1AmOLatncV5fVOuSeZ9EkWeTe3b412L/snHZn7kCC/6rJMTVP9VR7bHDxv/0xKDD9JSPYL1+2a
OYJ1nbPRh6Ea9eMqfs80DueCoL8+ktarJODqhI4WbXXQsLk+nwqYZFk5GSa2gMH1VcY26uBPRZbo
vahwzewogZM7pgcICxdXfpbSu0z2nuGj9yB4UJZoLxmLn0DB47Kw4+Pni2TJXoDOhaE5y9YRd6qj
LZHs+gWCEeCKGwaccK/BA4Y6IpuJotlZDNrx5QMNjongqfYm2sETY0ITiGeU1AuXgP8RnKc+Rg6a
W4ePMAANn5V3m+pCavQit9jq2zlArHPMbamdz0PMWOdnhxpk2aV7PI/FaJvBrMDtFBORb+iWHDW1
jVXNvtcsi7iYmwmaWo7H/DvWDyGEG3wHQyGC8IxU5dsE1iSI5xtcLvSuDIJ8vcMjGwttsaU44D0P
c7/0wDrTh2p3n8fAUzeGHuv08RILdKC0e3wkQnhxxliTN9JfD22FkWRtqe8vYUMPtM33e0ZW93op
3/pQ/trVz2smAS62ojGzg33IJiIdW3FDaI6mpHfVi8gTMm8dky4UW7UQXTeNWi4bTANqUMO5/6L4
CFYuNeFpSyPRudKYw1xsj2g/HPl8enHh8z0km/eNRHVh+K7oTJP8u63oEWbNaq9gGR6JdAbcD0uP
zrL2eG5v/YifBR00u/gsSEtQYedSjIVZsNqwggWMJoPl5OdKALNcpBVsnlM5vdWqeYOaST2BIdkx
DdAXSqtgxFfQe8PDNuGRXsNi5PrwqiESgNx/sWFwsKYiqUe/i7A+6GbPgyqqzmGbOLFpqXNmRaas
E0fP2xqKKzAdk2lrZzsLINVHHTWQQNoZf9REfc42ddE4mN2cwukhGugFed0apZ0mTR3xGqR+LA8g
0/lSOHNBeeIYzyXreDtnEFDfV4boUbzjS2MxEY3xWaA8EJLIXqsqmdbOR8P8+xQsjpiHYd6KyFTd
Bw5DzNrMqIroiKEmeOI/93mkXGg84gcPUr/DASJ3c20cKiaKVCIJjUj7MI1bKYtwtvAAq8JRkb/n
9laL1fVbCYGxygm5Z3HQJXZnel4sI/Ffmda7eXCzVB4kX3nBuseBAaV+0livBFyh49Dc2wRrTRlp
rH0mKrZnhD2P2IFwXzGJ4qP924YWqImkxgZmKsX0f+MxiL4Yc2a3+mFr3TTJiFZN1bcpr18YDy8c
Toam5+v22tvFlV6m/6/5F1jcBaFIgd+XOZyHmReVNS/piqLJbPLdPvldspF/eKXPJUn0jU6YmKVQ
zQfyV27ECnMWYb3rvHa1B/5ggo39DcdtBxfrAo4i0M1AKudevYCcRRbNlOcK2qX5IiZR9AIWXUZc
CXZOmq/R/2WW+jvGSEAkq2BFZz8VE7Weclh0osr5igFBnVt0whf9NIM6vNsSG0JmRkKE2BoJ7BCA
y4qt0H9muDHnzTUDfpxWbfvoBjdKfDqd0s9NKhIdiXbDUBSEsRijfB+CxekNTmxFuIc1cpjWvdRS
4r49SdIvA9g70ZLnLxbSPUTo0qlF1UgBXi8Ozjq0T46Do7IFY8TogFE7ofHr6Fo2BmK9gw3ANro1
YWbD9rdTHboaOA/jsBReMe9rc0qn0wsTSICJYF1IgQ77bQrOT35Crcss7NnE8uHoUSLUmX2nYdCO
Z0D9YAA8GQI283iaSRXWn4esqcU6+dvLPdFGxDMQrsDN0IgtCIca0zS/H65+M7nGp/28PWebsOPf
/lTCVf8b4PG+OflIQP5Sm/Ho3kPctSwK5V4Pm+jf1YY1dO82sSsDtfTCiVjt+eOkjRC4qnKa4yEy
lYCIE9Hxr9KEWO8dgtAdewAIKv2ikfPF2hR8ACiP1fswALuoP/Ue90isf8PgpRn/MGBUcuKY5aKk
6WaO3flWOaSqzt5Jn9pEuuguyeu2qJAWIkaoy8gj3NX7nSc6jQvt8ymZIVCsQ7wj6mlEW6Ps2k+C
katPh1ef0krW5mdq3qJYniUN3HEtQMEA2neQhQr1Div6trVwQtOI6kKTNE1tWHl/RhNnXWmG8Dp3
tjAFYRhy+saw743EepbWOG2Gxtq0sfOkqgSsKKikFKTkvtAOeJaYHmY7tBRebN2memtLOVsBbKUz
zAC5qOF5kJbiV875WiCGiQPNbXqcmIqOfneEDY0KDWeDWoIf9D5I1uCTEMrt2S4UKwrQeLzM3JlQ
Mr6XbqoaSfl6Uo0Z+8VS2Jn+/gAup/Cn7wikduGqOU7D/x9ksYtbf6lyvKhtoyqyoB+i1tH1edPL
cjSgIPiNLkE0WBBDEQJ0atXiB8Mvb8k+7jWD+vgmaxXOW0U1MYhIrBFvLZyt+IOIKhapsk/nQ26a
c8A8K8LMgPWvh5PyNGJifbHJRLLWWBSy4RakhZJExw9TuB8pjEy0CXNvjVoj9eVuqFF+UJ2BE7RY
1xjGUZCNLDhLXuCxZz2v5dY1pHt2CUZPb63esVAr0J9yP+o7vSClcSaID6+yM6A7IwL5rd0B7eWL
DGjK6qbk0m4UVdHDjL7awSLld7Du35jnGaLp2MRyLuWTBZWF7tXyBq19KQw+biYh/pj1telfsEAg
YffQWD5ze5K4vtEFyM2/dcO8kxxflfNXxPEph5xoz1jAosscZvzOcw91hi6bp9uTRtKII9rcVrGl
ZlDevUCojwlGVd3mx4kXSGolaLQaoBFa/PMCRsna1t8FEAcCW8VNwvbsc35BlxEYprSaorc8UZdz
mFBCb2ZPlLflLdc+CMcVxM6NQKRLicHIbf2AKAEw4375+79tdMmPSax5iANGoAjp9h/a+c/rsntm
zxnZE0avqwJTasqcVBuVqqun+JyghEY/5s2T2rdyPz/FVPHxFt4kyLUwESWuhWzP7t5IKJ6hvZ6u
EFYFsfPtgU/wonBvuasmv+qZmeTnuRZ0iGwuLplzAx9B6RSx7/02ZmBAtg7LhwTg4JLvxw8n3e1c
0H+Ck7yPjSb7hRrhX+oXyMVDhF3yfE4U7uf1+0DKun+mdiLfwDrVXfZ7EEmWN9W1kpIRxcylHTVH
fEDefJkTKATSbTRQvd94DCqq+YYcnna0s6UoSrNB8Kq58oaG58I2F/SjLNhIyoDFaydfzfV2S6Ul
qu8omKMCTEhMZhQrQrdUf14kASJ92VyDgje1lz3lNLUX9fz5tFNUwZXkzT0+mGHmbtIPq1ZWN5pk
8SIZdRXtbfYLjixLKXlxvBYGpqCbHpOY4hJ4nmJfU4xmdgE1TEEDuyTK2IPfB8m8UNNq60eC9ydL
mdB/E54jtduKdAATNMwhX+ONTXhtTLwb3lgc4VDOj7EbfsXHMJrSpyRjVY2UPLc1PRyaab8/+lPm
E1aXcuEcVPIiM4n3Ckcw2PQw7vHmAzWawhqZQB4ly5gIjFaRaIetFLW32scBm2PU0MYdVm/cUg54
+MSqp+XyAcIDPwYvaQ/mBieYuGnT7TFxyRoVIYMQy8S2pW/4Zun2FdR3mQBu4+f7D8JUo0oPKycI
xah7LQkYl8hUjI/gIYtFmNknM+rKssZKMaZzb8fDVaPxDv6OVcSQT1skXCee1FdwKDdddyar3ZXV
Do9xxUgVWepsu/ck5Sj075r2Lhgwo9teNbzwf5drvuJiUW0Otk/PsUI+8hKB6mM28oSY3mZX6O0F
ssKMY0RVAhvLdcqfrmgxlon9MnNpN3NmEBC01pq1P16dRN0J7PQhuYXMpWfTLZcsWSd5ZPZ1p/nc
spxZBSo3lGkOhJDfL+eenQjSKD8c6yyXQ4suohV+LtND7+qE6F7jsVPfAI0MOAkD0zxcMnZe7oGm
ICgRrp/QO4q8aS2mCE7jvhWAS32C43aSUhJUB/+H7qdE54NVzhF8UEurd51oEWMQ/IqNVM35hU9K
yeG3qXbH3h2isQKxH9mPDammkqG3l85jUgVuwPDeMiDPDhADMjI7IqusU/r27+Fy2RekJqiWdQH7
1HLP6JjdWmyULSMXazSdho+YNuDY2OJ10t4P1umBWsFmrBWoR81tO70pJZJQvRxfqfjKo1hFt6Qm
vu+NsF6oRAKiNM3TsTF1TmgDlcQzo/uK33JF0+Qk0hU2NNOM5DsI0cawqFmXi6emtn7FmlmT5TtO
sx0Hh+jvbj/Rd7b32LcDUsvvbJWyIyilNhVPwH4Agxk/chg67670PM9BkVrZjCOzsiQFrbW6m5RS
4dhTB7ZY2XDm6mHrkWaNqiBxXfF26+p/GMLNEa1w/Jc6GjoiErnWWvKWxm2wf1kSZkkFQmZII4wo
dExYYuh+KTmmrPTxVOjI7eQjv8IbcKLrQsixgvhFOUR27yuQexwRbus9XS6RqI8qP98ksM/0XQzV
kVX8A3xTcaiwaF8QSlPtFy7FKr17/mLUE0GVLSabYwtBUs4Ql/yFgu/Djb3HkMiuWXmD0MQiqnFE
Jpax7+CnnxC6atoOaWARql/sea+GQ8lOF+Z/0UoyOzIyqAeVsNiJyZSzjmFwzDe2+ZkUVKAuhDCF
3VGLwgYWjxywaFU8LMTGfaAR7601FDCqQwBwWs59NaHdFIdCQzt33969e6fZZQc7BjMLROBc50j4
pvvqrTsKn//aNRnQ0ny4nfTM904/HJwa3XZmDPD7FSnqiJJNKlLcXFCkYukbj7pm/0iNMMsi8hc7
yhjGhgh2tTBZX3Kmm9wF1v6uQiXhwstreUx+z630V2UwiYN6JmIhtjKMGB32YRpY87UQzZHsAXut
HMGTepcM8gtiLgr++xrraAlXL905zelQCBT0dA4m1e/inA6TFquNelUVYv4uGJeGTBjGx25x0R7I
/TbjAAM4kM+xdfap1HRh6PSomVqH19amTvalnnMCUSwKtkXsy7BexssZ/UiEuEz0QQW/WjCZNPYG
a8wxXtQrGWKDl48+s/lQ2oPAsINupSZ7SSJC0EX//ySka9pcLurWBb7wnIs7nwrWbtCa5RhRIEqA
Hgb3ZpQOfWoxoPZTkYMB0+EMEfcSgTVodLzi88cRmWo8hWUJZNyErYqCW3cN/sZyGeplAapxhOSq
XCwGvoI9KSUev+QtQweaAN8SU8420qCHLjlAvq23fh5mpKfQne+UwnaFrFGHUIcLpo8jtBTje9ZX
mLmLae7nF241Bmqu0Lx1QKoPZ5bH2abvCkAIN4JSGbLdTQOsY12fJdWlEOOLpXqSJqd0dqX9ArpU
7uKCHwJL3W2dCbhQh5sjdkhjrHOqlxM3xYgs42qCNCmUelW4siOvPzv4e45VimMTDuHbgLxfWRIq
YI5QAwpKcUBdaxu8x0L/Poj6r89c26R1dYIMl95UnX7qnFNK8H/gFxKupOozBujkJkOLkN0zk9fr
Y1MFVXxYi6P3pT2OH0B6TQfsvf6nY6cwGCgU+GRpO+x5w0alu52MjyZYYXYoLaUfhrJkIdo06OPj
tbpXDLar91R4RtQ7MwsWdBIGVY/0lIckptE3D9Zc9PtpPVqAEiT4PLlCCh6CxiAygomRU7vmJVFn
ZKnVXPHuV+Bj0F+yuaPNU8ZsC1fQf1TDaziQSsomdjV+i8QF5OCpAx76MxogEVTtJK21Cb5S0GTO
4uNn8XnWhjQ0W5qaJqRfAB+UPHdMSjgM9NxkiUSt/3gKJTiH8WAPEAvkq5Nll+OKl7He/5icz+P4
RqK+guISdpSgG7lu5Gf6XO9s78Ug9YXjatyMzjImgbsMjU5dj7vrfTEeeIkelO0yIZCRBTumGu8l
A/tfaR/AwYf0+WBliaGppcZfoKY6rHWQ+45oDHHdZnoaLpA+9eS5pRTUxX1R0O0X/ofK51g+if/6
b6mLx/CHa5PGuU+fuc/V57F4gRTsVAWOkWLyEl0bNyQL4cFwEMlt1WqoGlvbyalXAxnlTuXBPah6
3nMo9af6s03c/a1rblUAAiExeiVvgxhngPZj7WK/B/60jzhnWa5o2ZAql+WrnbYvgCi3dJsekH07
akqPAi2clQ7fn8HC8mjy3OHsmV/olqmuhgoX/kHorFDv3VbQgsu41W67mBcE5L7KkOsvSRjYs+eH
58uACEsHLBTg0x/EwCkjfkmcImpHryx5nitjBDlQMUuQ6dnP2jPSk9YR3uVuwmFbB1PwjZIjaWEN
TaMnhSprfnw8Cjb+PoK+ZW+HlgedC9NezB5uFhAZBAEmo+iKF6Mj+sMJNaJ5q6SLI1HNwQI2Aykl
ryU6d4IMaJuYNG2mwYbAWUbsgQxv0H6n7wLTntp2qsEzqlMzvwU0r6Xi0LB4gRGP+H1OzJRi5AC+
gC/To5bIckgedgNr3O08UTDrn2l8SKd2xeOjcuOLroTYHj6vzETqvOBG/IF+nf3e4yWIdKuErk1e
b2JzZtomTzS6xmQWkZmJcU/BH+xwMgixOp/N6CWZgabnRoCbo9dedre8xZTYzoFOnw9ldQRucWH4
1iSUwj4raaR1q6wIIKZC1j0DoWYq0ttHkf1aJViSOM4n0ql7+oi24PelTXJiEaHPGokdbgjccpx7
xTWDxppV18CzSCgcvUvksuGA8Hk5AismSpgOXp00mSwHHAVF/mTo8nZ5dMCK2DTYnydA5RpiypbI
jo2I2NP0GtolBAfBtUpEyhyEmA3rEqx6QJZJ6hYVBmVrHf1N3AfMXdxrcj4tiCW9oQtM6KvFXQPP
KNe5ns56Bc9S40keIvBOSv5lIujj4N3G7GTvX3/twC4Ilm1ayh5poKqfh3rJ4kQa8Uts7WvkCK69
GgBhT+FbecngxXNJ66u3khxbNt0BYK83ACAhwe/R3lhUVmd2D5XTpMIZSyA9V5LETh51ZM7+nm5l
AJuOc2vo8VpPfGardmbtVbhtbIDDodQWByD2lhqkZ1KcG9fVa/nU7OS8mPq+opIMZXPKXA2k9ghg
RMyKwLLvKJGVHHM0AfpoNMYkFfnYxQFx6hmcOC3lfza+GAsmkQ3X9VB3IVd+S8TnaLrbHGd5cPWa
r9dOE+bM7jeOH13FjsLCGTngZU8IuLHZylrcjTb7RCjZV5uDVo+30++dbNFnTIxHnwrnXqWyqsi9
kFDiZAWRAa57xzGB84AWAHtrtxB9lRPWhTJCEdWYC9SWre4Xc7DAZQ6pRVy6KK/+EZ1O7HZiVwB8
uhaVZ5tzDukIVTCKnlK/sRdKvFyzUVYXqWRH+gd2mvtCrjjTtI6YtbhLK4jAjDAwEMvbZypT7iyw
QUdTOTbq+fbi/47V1FfdicLHr1ynbQPQXeONaSWaIl2fontTXbh0uJDlDPAqOZjSQqndjUpSIseJ
tKFgPYPBD/p8sSGL3dXU1muqM+vhsTJkPuXDmkfO9085TOhX9fmzH2HXeGnNxPNFDisC0t8mJ7EX
zztzJXHzYfqg0qy/SdrPm1L+7OSYIKjnDxUJTfO5lKWdccFdi0iKT51jxSpehKtUtEt7CgEUWbaf
b1dXbTptxbJAvCOqWOBa8qrgKxdTLzw7yVKfoZxevDnMcoNFCxYRE9j1jlwB0GEYok3Z/6gnKoBy
hr8ch8jwq2pq1IT2Jf9/GkF47G/RVwRXdmdkVWQkffR46OlPQ8HH+U7/h4XjwCcJQE/jPrmIsF11
W7qy/h6OMz+kHWpyo7b1stMoQyzP2HEZN/OiceZOUKQzMvWkRt29UjxbpK1Qj72CwVpUSA3XWUkK
tYbI9+Pdckj10dPlmtavgVMo/mFCmWXH4pLhwQnh+3Bfsym8014Kd7uZpJMdohsxtRRIs3Zwxz2a
JCievnOcuFyZ8p2AX7iJwGC0tR/+i6t+giJp/qorf+48S3KkStoFcf71Sdrr6mitEppW8H1rHRJ9
p7qi45qAGHX5nY+8IdYPe9JmgIbih2NdS9c2c1DC5wPJBs71Th4V0vjdnXt0IkPiBbQSCpur/8tG
wlAKKAM9DZsyJsrPugjXIvMv3x1pB1TXu9Ls0hSuQ7WEootcI6TYdRt0Ez2iIzouz7d9MbbdAeQh
tdnrW5qf5brp3Nim2hqrFjW45wMNMVK3+7HA8YceHTOGpL7u/H5q2wSvIyWlEEaZEF7OIaGDE+/g
WTCyMkKrUMKUSbCY1KyTzBzz0dTWAPr/osR3B1aZ9/0D7rT9GS90R1S6IwkhdzTkjHYThpw0wnAL
lokXKlhYAkKovgBU9hRMO1FWJ0KRBurFRwDW+dbIQRr+H9L18AT1NL9urWJ8M2+f8klZMr80hjoB
R6TaJMXve+h60RWQrZPpRWLGNrG+rHphC4rhKSlnKwToqV1SLSI0Vgjmx3tyY7g8RmTA0ita2s+d
rAR3w4rrw3iLE2lGydY3zrJ/vjhXAxdEBHpoGUR+7deWfwYne0ZsPOTFDYcg21hUWcm87/I5bnJK
hUh+7iL1RMRq13va3E6ZLWnYXlYG941OmHKVskYloACCfH7TD5gRWYB9gDMrcxjnxXo/lNB95a4N
B0dGWm7FkIVYiOr4Gy1uB8zabFBebLJajsAbAOwg2QOZzxpPOnd6bujfj1ycpd9/NMUiBxhPYk4h
mjRYkgm8xzY/8pjFnZUX2uPae0sDqVnzXsSLD585FCF1upquMYTXeJX6jgvSDiwwSH9IaFSDzxO/
XWbm2JOHN1h/RvLnVIQxrWu1qVufykdk24BZo5FFvSiOqRh2oaxrmrMs8G3LUP9Xut+Fi0EiLaX0
puRdu+BP7qdJnZFdZ1FtalEcVc+K6Rxxkx7L+GwBaW4vIa/G7NjBLytO83LfhJTVA5oc+PrSSaSt
N3XSnqUI4EUf4DibblUKQZgOqMpwlWdD2EKcSRBCtzbTjrThxS1d+XTI49ERSUF068HXcfTDtMUd
KU9KXN3YB8GP0VfTazvfqqwYij4RbRFGnh33U/WXPXCuzXQTzaTwqvew/S0VqN4P6tR3DUbI9xAu
b6paI5oWhpo8g/EzzkdJnwAs1zOSSgl57Y3qjINsxmavXR0tDghcKNugzLnPozhtDav48i/8jEne
npXWSCubRk3wF2NPZKqBnvz4DGubHqa+SfToToYLkkMxwX7+Yv34TL1WC3KJmWTmYDULCCCYAcFs
eViWIEnasZ1LusFnAdnG/chxR6qLTcfdlcH0d7InaNbPq0sCTj7gbfpqXGOgu0ZFAWC6/z1mQAjX
B3KEXrkY64Cy1xVCcAmlHCtCjd7+UMOe206JgCJxdwhJitn8r7hvpeaqoCTq4XV1dJhoLQFtdZZL
wY/IjdjRysZI+kRYwOa6MUf+FqFo9/bZ2xTLaA5cvibWsJdA8ce32H9hqyKeCjmY6V9eM0yTZ3YT
dX2nbmYu+y9BHc8Ap4WDiEfG1P0i0pFFFRfIZ2eoQxLlV2Y3MKH8sru27BrpHvlIxU8t4ESXhn48
heUDb/aJWn24TI5M7YdFtcn/Zy7oDLQWw44uO1zRhjZlLMQpdK61HBspGsHwoh6rRZCI2+DzDxhc
A6x+UqjCSuJCF69IcKoHWe23DEYlMQpxeMEi0QAmW3pSBIivuTj+2glDIXBaKc763TxGOZOsnkWV
qSva0/6HOUXOdiCbAV7jcWorqypMWia+b15e7Q7fkM2Cc56EzPtRgJcHL8GtNKu2ew/NXJCm8MlZ
rtqR+I07TReM8MbQfCocoGgTaZ1HfxqEhFmVh9Sl5saVnGVCfqcAjN7NgNqqgl4NouENwtgy42xM
v5uoQar4KO7iZll+6zTwUIvbAexBlcr1V4lNKrQTBGTOWtsj1ecLZwOk56DwSaM/aS3USVwsap2L
7b0oW386Ueh1FEHNu4gE12JqbqZlKRYMseVctK07wKn2dm6bNCi2vIt+Otvepl2URr9HvrZy9hz0
9vCeNy0sg+gU1PYVWI28Fi/7i6Fx6OuXBg672wuM6o7PXIbLZEUhB8rpyozRQ9abBSMnz/MTe2bQ
7mhydcfXN/1K/8CfXwlPRVVfZkAp+0knIKAQCZmQmINYhix95QoX3pYCDdhk5oRnPuA9Qgy9Uh6I
u92ZJGiIWyIgFFOklbjxscYf0GiNpe7vUWUgbIuCAkhpHxXhwu+bP9NAnjQOctQtiShpJ/+C+Tiy
XrkgK1FNZWFamyQ5IRbCIHnVubd8HFFXgIN0LR4WxjVQkkwoqN2k36RREfBOVZFM7WVh1cHuNcJ8
GIT8li2nLOgRRGmhXM4kRgNqUgbCPowTABetYPdtw4jf9EOvd+VEVXCg+aVi/8qcCtuswVT4h4jl
ckjrapddOWnEZah6mkwbZulB3vGvV2YC0oMS37kTlThcwiAgcY9Dp37q8RFzzAo7XN8ITaHab7hb
zrRIUzacMiCznR9St+Em6rLqSFCgCC/MEt5AdLbLdykAD0lwXW9RZ6Rfn/RVjtADsrmEajHSfYHH
HGAQ9nnDJimLEeDSJFEKu19LjxEp7Dn85qScSVrFFIuMC+d9aRC4ZPvUVk2MBwNH01xrdfNXF535
mWvg2LeTDQmtqdNqZ8Omdqcd8wEL/K7jTY/AdgLLfkeY4Shep4RmnEtovfua6liIZIT+cfReopuj
OzHnievbhNBkvRgbHvvTex3J9LDyH514i/NlUiuiciAGQx67WBXYl5yp43mIc+adJSaL440CGDJs
dRzsNcIeMEwj1a2vOVS+/VQykgZ5YBDng3/N9iVxidOuLve25w377m3ytXe8l/mgWu9nilpHwKvc
uxCWAUkYjSrwqXisNJYVWia4l2yrPscAp9cUVJ1lRn81cSYv84kKmHLgYWjmYDDNEfozBRMXe6wU
/ehN8bDnbUKISZqK+wQ36V9+Fn0ltc+AYUMHYGFLnZBs3PXDyGonvxbKV4gNzE5sS+0ugLsA7Bxn
ePqO1dMvWxSFpM5g10yPu0OjGu367XtnyqHY6xtEnDg3HWq0IraVSB4tk4mZ15z57iEQNV8RNT3U
E6NEtfVqJDve1HwXpOOX+GVkPUXXPNLk+RsvFwYWQqNCWrkwFE2skK3GbakWSrSjSJgX+LseYKPo
VgwLaRvWG4s7rpT3TSCH9qjQ3HiT3Go2KSIwt6ZddvIpFM5ity0amaEW8xfKzEZEtoZ6tgxlGrtd
SSNnz7qwytH40flcm80aAKPEyPFQMUAODsJMCb7BtoenQ9IaWP5mhACUP8pk0Hf82eDMFeVzPWcm
EYVok6MQKU/KX6FiS8DuWcZ5Im1wbU8QeZKPhEE8Ro/ZjWx0d+6Xpoqg0U3uXUvYhmGtJ/8Xy4ru
jLtHDKDtIJjiRqumtXC3+rmlVWHRwkw7Q1b9alR/QWtEEf3gqnWmZHrJLXNSQmyrtw8OVywYlF50
NSBrUyKxHf7XVMjUo+iOLNh0zgK/PX+io693rMQ8yYBCRpKxopNchjb6FKmU9Vl3gcAOH91TZPoq
Ky1d7XQMCq9FryL9rUegXHqFCE+dMnYqmfuMF8suRzeKIWIAV7ryJcBQ7duGxxwnZ3Xjf2+tUOD2
hrVG1NcdysFumg3RnaXuckhF3GHT2ZoV+enWIeNhXmyVS4q/slq4DS8kOCwxMefwjsHXtnDMrZMm
wm64GDq6fu0MPiPPWkht6QFRhj6WMDzNX8wXVhAFFvVvOvF318spH2aYMoBzZ5NrMFn2NgeiZ3Xe
NbraUEX8vuo7ziGCudPlhynaGAz3QQuolxdeWq/XGkQMRIrl6v9O8wWdwew9BHflDuxM1i8e+N+o
z/LDhXODhz3STf3UdzMPTQf5Vst0wvPZmMjVpQhhGnld4h0MfgVvP0pEDsh/jRAiT17ACiJdBhf2
nDtAarEf/ecZEzMxUAJ8NBi7STDIoidYkKnDa4U8z7ccIYo1gDhkQfj4sM1jKXRR5XVWMbw88Fxe
tfpCPV73hQzpLLsSQrynV1F3Ja6qlEbhbsDG6IkIpGNO8b2LY5vEUJIuh3d3I1kG2M6gs0yO6l/W
CEsnahh4JybQTilyj0pq65h4EqX9Dw4tYSMv5FYvFpo045jsQiUjNyQuI/3LNTKLgPqihcdlmdNn
K8MpRxJ5nkbZH+swGwCPu54bZmXZOtiJ7Ek3PFNZBGTyoFEmEgriCBsijEDIO6LdhSdH5NSHe1cC
rQ23DL2Dal4qxRqgQ7KbtmK3uZ8+epeFQsJ1X73foYkUJ1NXBNe2o+lHTIxHecKvkfy2yiUvW9KQ
ZoVDxyK1UbyNBzB8c74LdpwWjyxBtk/nxiT0n+KUF+Bja+fnN7ff/DxCTKgNrA7TOuCplY7bPDfT
oG4L13M1Tp0AMGLW4G7P7+BbfZiFKh3e+8a94t/LK9TbVa5MnEDdvXrNtKgPr9AbmEd6XiBfDr6F
Ci3Gu1XHllTWIVCn5Q4trPxXSs9KY5H7nEvyv85Egie4grKZdqcmZbhlc/xWn89rfuzScbScwug8
JfdCCEclLNB0Jqbv5IhYj233YmQoyHYfVUKAvhFsNkoduMFtzfRbtNgWZMdVXN8ZTIdXg+a9fy68
JcgWS2ZvSczswNXAhEzF42D60jWsk7taNJeLnl6I20VibR44OgFFQOu7kKa2ZW/VvE93FpIgNWXe
9X3+DYsA36vbiggnKZWJXlGPsT2w2bdSB/tVxv+9i54w02V+P0eT6wlX4gQGf+0toLSgXlK2t9FU
BU2iFR5DY5fkVjMIMX0rFzV7mBbbBAKFwHCjHZNWCZQF/Nr20DvM8hY6OwSh7DVmSmEKCgWOcSUY
JMcYWBb5auhIKLyq0h+zBNtAZDvzh+j2YFBrkT0D8rZ5+uy7xG4IOX5pHYvcN81qXQOlSUgiMAyG
y9cin9hkNSJGCaLaulTwCAydvAgdTWOQQwenqPSX/a5HuQUzKcisCTOtgXKGAQtJa8bVa2H0ErQL
d69fA4uRvsgNX7RDlhQuiYLYZGCiLr+7JaOMGmOfF/m0RNNJYt2WFkFni7ljiENJ/5+25ppx0WN2
Gx489qThfzLNeGLOiUzax8Z0P+EZa3eLhV2PY06Ag5bLJwEtO3wd74mbgcGswck3afo3ixnzYXDI
m+14HTlI+ugscnVoe56fqA6mHy8hobJj7UaJ6Y1HJC1248nA4gpDmxCndsl1jQFXsX2rfaI6W79Y
MCBlIlXHGi1ut3y/0qGUWl9ZCo7c+a1bYvARitEgeYxVbszScySOCaCXNQCaW4ColaSJyKyeF8ys
8sISUTLGo0U+HLQ3spkuIlkmMlHNEuD7ydnudrqVrpvcIhfdzDPaQyBFYBWSXgcwwbvSggxK41cQ
GjpZHBhdtYWSmJ4EgaOV61i7Ozw/ICAU1o1593DWEySa7QzyC11Dqegnzbj3CDgEereeDtQocQM+
kuZpFgy0Bf5PeQYE1Rbt5W0V0wko4p+ZtYaSZWS2KOL+AfP4LE5mvu1cd0XkXOKEwYkSdAs94K30
x/uswGZAfUB3ISYqbrMauJap7WV5D35TC73jMUXLjzIRZfaCscTtQxKjUk3zMnP8Dh136PVfKGUY
88rdeUfrWWN/0qMqiOHrb0pB/EzePvsPtavd21NVz+8PX61+s1RYp8pAakkXhMy5YfvgCiHFrxLI
Ndmot3WWGcNSmmNgQ3m0KQ0qbGK8ld1F9Xj+TD4rgkuV9UYVN3aZQ2/g186+MeAp5usYe48U2tDY
YY7actevyji2cp7ryE3/xEONEKRFGYNe16Rgk/2eXiuB3tmfmECrK/v+H0E1/vWHGngFlu0EbL/z
FU4ctY/Djel2SIYPFa/RgC2O9q+k1f8+syGL185B9sVocU46l5DRUVnD3OeYGgZNpDUxxFeHbnBU
U8jfp4NrJHi4QIKHO+KiUGeC6csG/2VIDv/8D28NITzxA7nTl6PvnSQKgwJFVN9vtu8iBy7RN0SN
dWM9tvIETCwCQrXJf9tDIFfK5Y93Xu0nMFGIQtheUckJe1qTbb5nPkTZgJD9ur+lh0aRVTWwdjaz
yYN4q3/DN92o0sIX+5ZIh0gIMgM5m5lru1OqrrQ/dRxx+Fljub0g0ryzgIEs+SoeH3E05P0hFK71
0h/2y/mROU2HNFQIXhuSH5muWM4gYChxe46wzuOTiU/UPrNf9uJ3w5Gu//sMjks9LobmTdxQp5x8
B7hV5SRScoQrnuujsCheJAG0k1H7bWqwCTkbn+XgzUnEg7GWMIXJV888E+sPEkikpOCcFH7eb3xx
ajbKWRGgk7kK7t720ESGTg89H88lroCi4K8ch1zTZ2jL5QJ/VYEF1HPc62p5FNXAhnpfRILdS6F8
8mLpIDP9aMjkiDoas67PvuYJZzSTcq2AJMlZod++wh/919Nad/1NrsR+3DvseEOCjsVsO9CDPrTS
3Uzo3hK0mvMLdUxErWazQ3qaJGOJQ4nZVPJrLyN76ywDENEFbawUprqHzRmlxHGG/OehPLDyLgib
W3+B6GLrlnI9BazMaOGzJvk5Z2b9vKixQxB6wKshLLb8WfNXKEfqyLJImL/sJ485tPON5zXaYC4Q
Rf8uttheSfGPd3conUwja84+su3ZEw5kzn51WpfKour2wg/oU5kWZ5MD9d/0RE5Z5ZA3Mw9br4TO
q7xQu4Yn2WHBVrs+ILcP3wBtGXkc3p+Yao4ZZCTFDJ42HYuYgg6Y8n5q6zTy0WbzvQ5N1v7DwRF+
SM54iqJWnKNCuDS/K+Vtay5UBa/oZJ6NNKsKFYSiMJ5jjDwVg9fE/SmGUrRIAcBIseGOj3YA4VJX
lsguGKuZ1L9Qc/XAWeE8gw6Q329jN43DoORQNp1dXKNqB/1tz9mXAqMWiABtKfBtrnyxlPFF7mMU
iA9llWLYdbQdjsdmR2tfhHBVbIzUL5UHxmXaZCLCIeZhS5PPC2/sD3vJNtbJlEJb0NBJXYC5iner
kH8wdfKjNFHR+jnd1t/nZX0rk6+XjDhF+U01JG0IqbxZvTygNQXWZ+kHh2xl6NLEppmeAC6y6tjh
M3m+EwRvpbXcRy//JblM1qS2xLL7igm2vD+EkMOAWDOVb40ppAJVL4myq0pwhjSvVXAFQJZPz/ei
vC/0kurpu/Avb0Tq9cHcx6bVtgKXxFPHseDB6Q6+mcyKyAsmG4N2Vowxo4s98YdES9fZ8LPuZGP/
TO/i7Z930Xbfw6QejfrJcuhCzdz/4vVoVNJigYTJMyCKzH4ojN44tIMlsa860CTmTxh0DuLX5WyB
GpjrsAIxJIIj3T+60XYu07D5BtkSMcqslrtjyv8No5C0FHNma0y+m0ztOODfYjElg+4ZzRLmQDAY
A7Nxz8s7chvItlEFzzgbBEacCPY3V/YNu6EcpPFdyAMCvZ04VndWS2f9a5dWyuB4d3g2p/4CrGk3
j6HG9Rp6FP2fIcr5YHy98MmnLZZmqJ23C5pffUwQGjJaSm6Voii3IoLUsXYFWmzRL/PKQyAft/iw
W8OBIAmhAFndr0qHtno1LikBEiaGLLgESB/ktH9X4JjpPW16Zjmw17XmBTohubsCivjz8fmPhksh
RKT1kxloCBLAZa1vguhw7i7xn8Nm4JjP71h/JJ1yLJIb2I2CepOyiDy6E3OtJTSukRphh7Q7uqpT
GAy6go9+iz9HDGfUTbWbYWpDLmUhNgFNRC7LrIr8wtSYupv8vyPRzxhJcWKxZoAHYfSL4ger27uI
v7wEAou2iHqCy4iS7i9yGHkriQu8piKhjNdY+Z25yQ91ZYHSLI/sNn3LYXzerXoC6SZsDwA63Wjb
mHofQlWJsUU4Hu4EOJ5OcZtIVH9qwSQKdYe2K53Dqt47LH6KpmM5hl+qAgG+1C1vIDoM7KKeEo/0
CO73uXi+9zDMPGCLBM0AKA0NNVo/WJAsTO8yAIUQbfuchAyGrdOi3GtBFFel9A46sp6fRKeEibjF
iMyYrLpkow8xGp0EjVfQlIIbSOK+R2zIeeavL6COCPjKHHYtjQ==
`protect end_protected
